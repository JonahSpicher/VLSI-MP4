* SPICE3 file created from branchl.ext - technology: sky130A


* Top level circuit branchl

X0 a_2390_n90# a_2370_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=1.5925e+13p ps=7.77e+07u w=3.15e+06u l=300000u
X1 a_4700_720# a_3710_n90# VN VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=0p ps=0u w=1.4e+06u l=500000u
X2 a_n250_n90# a_n270_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X3 VN b5in a_6330_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X4 VP b6in a_7650_650# VP sky130_fd_pr__pfet_01v8 ad=1.1025e+13p pd=5.11e+07u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X5 a_2060_720# a_1070_n90# VN VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=0p ps=0u w=1.4e+06u l=500000u
X6 a_7670_n90# a_7650_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=1.1025e+13p ps=5.11e+07u w=3.15e+06u l=300000u
X7 VN b3in a_3690_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X8 a_3710_n90# b3in Vbn VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=1.1025e+13p ps=5.11e+07u w=3.15e+06u l=300000u
X9 a_8660_720# Vc branch6 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X10 a_6350_n90# a_6330_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X11 VP b5in a_6330_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X12 a_n250_n90# b0in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X13 VN b2in a_2370_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X14 a_740_720# Vc branch0 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X15 a_3710_n90# a_3690_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X16 a_2390_n90# b2in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X17 a_6350_n90# a_6330_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X18 a_8660_720# a_7670_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X19 a_7340_720# Vc branch5 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X20 a_5030_n90# a_5010_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X21 VP b4in a_5010_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X22 VP b2in a_2370_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X23 a_740_720# a_n250_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X24 VN b1in a_1050_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X25 a_2390_n90# a_2370_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X26 a_1070_n90# b1in Vbn VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X27 a_5030_n90# a_5010_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X28 a_7340_720# a_6350_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X29 a_n250_n90# a_n270_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X30 VP b3in a_3690_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X31 a_3380_720# Vc branch2 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X32 VP b1in a_1050_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X33 a_1070_n90# a_1050_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X34 a_3710_n90# a_3690_650# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X35 a_6350_n90# b5in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X36 a_1070_n90# a_1050_650# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X37 a_3380_720# a_2390_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X38 VN b0in a_n270_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X39 a_6020_720# Vc branch4 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X40 VN b4in a_5010_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X41 VP b0in a_n270_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X42 a_6020_720# a_5030_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X43 a_4700_720# Vc branch3 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X44 a_7670_n90# b6in Vbn VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X45 VN b6in a_7650_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X46 a_7670_n90# a_7650_650# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X47 a_2060_720# Vc branch1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X48 a_5030_n90# b4in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
.end

