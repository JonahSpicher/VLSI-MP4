magic
tech sky130A
timestamp 1618370474
<< poly >>
rect 1920 -440 2060 -95
rect 2020 -460 2030 -440
rect 2050 -460 2060 -440
rect 2020 -470 2060 -460
<< polycont >>
rect 2030 -460 2050 -440
<< locali >>
rect 2295 1170 2350 1305
rect -805 1060 -250 1120
rect -310 915 -250 1060
rect -2245 790 -2160 810
rect -750 805 -695 825
rect -2245 -385 -2235 -365
rect -730 -385 -695 805
rect -310 555 75 915
rect 250 -120 295 -110
rect 250 -140 255 -120
rect 290 -140 295 -120
rect 250 -150 295 -140
rect 520 -120 565 -110
rect 520 -140 525 -120
rect 560 -140 565 -120
rect 520 -150 565 -140
rect 790 -120 835 -110
rect 790 -140 795 -120
rect 830 -140 835 -120
rect 790 -150 835 -140
rect 1060 -120 1105 -110
rect 1060 -140 1065 -120
rect 1100 -140 1105 -120
rect 1060 -150 1105 -140
rect 1330 -120 1375 -110
rect 1330 -140 1335 -120
rect 1370 -140 1375 -120
rect 1330 -150 1375 -140
rect 1600 -120 1645 -110
rect 1600 -140 1605 -120
rect 1640 -140 1645 -120
rect 1600 -150 1645 -140
rect 1895 -120 1940 -110
rect 1895 -140 1900 -120
rect 1935 -140 1940 -120
rect 1895 -150 1940 -140
rect -1925 -415 -1790 -405
rect -1925 -460 -1915 -415
rect -1800 -460 -1790 -415
rect -1925 -470 -1790 -460
rect 2020 -440 2060 -430
rect 2020 -460 2030 -440
rect 2050 -460 2060 -440
rect 2020 -505 2060 -460
<< viali >>
rect 255 -140 290 -120
rect 525 -140 560 -120
rect 795 -140 830 -120
rect 1065 -140 1100 -120
rect 1335 -140 1370 -120
rect 1605 -140 1640 -120
rect 1900 -140 1935 -120
rect -1915 -460 -1800 -415
<< metal1 >>
rect -2245 1725 -2150 1745
rect -1935 1725 -1680 1745
rect -1695 1685 -1680 1725
rect -2245 1100 -2145 1650
rect -1695 1625 -130 1685
rect -805 1140 -540 1205
rect -670 -180 -540 1140
rect -175 1190 -130 1625
rect -175 1165 5 1190
rect -175 1120 10 1165
rect -175 925 -65 1120
rect -1265 -215 -540 -180
rect 250 -120 295 -110
rect 250 -140 255 -120
rect 290 -140 295 -120
rect 250 -205 295 -140
rect -1925 -260 -540 -215
rect 100 -225 295 -205
rect 520 -120 565 -110
rect 520 -140 525 -120
rect 560 -140 565 -120
rect 100 -240 120 -225
rect 520 -240 565 -140
rect -520 -260 120 -240
rect 140 -260 565 -240
rect 790 -120 835 -110
rect 790 -140 795 -120
rect 830 -140 835 -120
rect 790 -150 835 -140
rect 1060 -120 1105 -110
rect 1060 -140 1065 -120
rect 1100 -140 1105 -120
rect -1925 -295 -1160 -260
rect -520 -275 -500 -260
rect 140 -275 160 -260
rect 790 -275 820 -150
rect 1060 -275 1105 -140
rect -1140 -295 -500 -275
rect -480 -295 160 -275
rect 180 -295 820 -275
rect 840 -295 1105 -275
rect 1330 -120 1375 -110
rect 1330 -140 1335 -120
rect 1370 -140 1375 -120
rect -1925 -415 -1790 -295
rect -1140 -310 -1120 -295
rect -480 -310 -460 -295
rect 180 -310 200 -295
rect 840 -310 860 -295
rect 1330 -310 1375 -140
rect -1760 -330 -1120 -310
rect -1100 -330 -460 -310
rect -440 -330 200 -310
rect 220 -330 860 -310
rect 880 -330 1375 -310
rect 1540 -120 1645 -110
rect 1540 -140 1605 -120
rect 1640 -140 1645 -120
rect 1540 -150 1645 -140
rect 1895 -120 2220 -110
rect 1895 -140 1900 -120
rect 1935 -140 2220 -120
rect 1895 -150 2220 -140
rect -1760 -340 -1740 -330
rect -1100 -340 -1080 -330
rect -440 -340 -420 -330
rect 220 -340 240 -330
rect 880 -340 900 -330
rect 1540 -340 1560 -150
rect 2200 -345 2220 -150
rect -1925 -460 -1915 -415
rect -1800 -460 -1790 -415
rect -1925 -470 -1790 -460
rect 2255 -890 2300 -50
rect 2245 -1020 2300 -890
use biasgen  biasgen_0
timestamp 1618201460
transform 1 0 -1545 0 1 1140
box -625 -565 800 605
use branchl  branchl_0
timestamp 1617823527
transform 1 0 -2035 0 1 -1155
box -210 -105 4385 820
use dacladder  dacladder_0
timestamp 1617750207
transform 1 0 -5 0 1 1655
box -75 -1780 2355 150
<< labels >>
rlabel locali -2245 800 -2245 800 7 Rbias
rlabel metal1 -2245 1375 -2245 1375 7 VN
rlabel metal1 -2245 1735 -2245 1735 7 VP
rlabel locali 2350 1240 2350 1240 3 Iout
<< end >>
