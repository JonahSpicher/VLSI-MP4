magic
tech sky130A
timestamp 1617750207
<< nmos >>
rect -25 -435 115 135
rect 165 -435 305 135
rect 355 -435 495 135
rect 625 -435 765 135
rect 895 -435 1035 135
rect 1165 -435 1305 135
rect 1435 -435 1575 135
rect 1705 -435 1845 135
rect 1895 -435 2035 135
rect 165 -1105 305 -535
rect 355 -1105 495 -535
rect 625 -1105 765 -535
rect 895 -1105 1035 -535
rect 1165 -1105 1305 -535
rect 1435 -1105 1575 -535
rect 1705 -1105 1845 -535
rect 1975 -1105 2115 -535
rect 2165 -1105 2305 -535
rect 115 -1740 255 -1170
rect 305 -1740 445 -1170
rect 575 -1740 715 -1170
rect 845 -1740 985 -1170
rect 1115 -1740 1255 -1170
rect 1385 -1740 1525 -1170
rect 1655 -1740 1795 -1170
rect 1925 -1740 2065 -1170
rect 2115 -1740 2255 -1170
<< ndiff >>
rect -75 115 -25 135
rect -75 -420 -60 115
rect -40 -420 -25 115
rect -75 -435 -25 -420
rect 115 115 165 135
rect 115 -420 130 115
rect 150 -420 165 115
rect 115 -435 165 -420
rect 305 115 355 135
rect 305 -420 320 115
rect 340 -420 355 115
rect 305 -435 355 -420
rect 495 115 545 135
rect 495 -420 510 115
rect 530 -420 545 115
rect 495 -435 545 -420
rect 575 115 625 135
rect 575 -420 590 115
rect 610 -420 625 115
rect 575 -435 625 -420
rect 765 115 815 135
rect 765 -420 780 115
rect 800 -420 815 115
rect 765 -435 815 -420
rect 845 115 895 135
rect 845 -420 860 115
rect 880 -420 895 115
rect 845 -435 895 -420
rect 1035 115 1085 135
rect 1035 -420 1050 115
rect 1070 -420 1085 115
rect 1035 -435 1085 -420
rect 1115 115 1165 135
rect 1115 -420 1130 115
rect 1150 -420 1165 115
rect 1115 -435 1165 -420
rect 1305 115 1355 135
rect 1305 -420 1320 115
rect 1340 -420 1355 115
rect 1305 -435 1355 -420
rect 1385 115 1435 135
rect 1385 -420 1400 115
rect 1420 -420 1435 115
rect 1385 -435 1435 -420
rect 1575 115 1625 135
rect 1575 -420 1590 115
rect 1610 -420 1625 115
rect 1575 -435 1625 -420
rect 1655 115 1705 135
rect 1655 -420 1670 115
rect 1690 -420 1705 115
rect 1655 -435 1705 -420
rect 1845 115 1895 135
rect 1845 -420 1860 115
rect 1880 -420 1895 115
rect 1845 -435 1895 -420
rect 2035 115 2085 135
rect 2035 -420 2050 115
rect 2070 -420 2085 115
rect 2035 -435 2085 -420
rect 120 -555 165 -535
rect 120 -1090 130 -555
rect 150 -1090 165 -555
rect 120 -1105 165 -1090
rect 305 -555 355 -535
rect 305 -1090 320 -555
rect 340 -1090 355 -555
rect 305 -1105 355 -1090
rect 495 -555 545 -535
rect 495 -1090 510 -555
rect 530 -1090 545 -555
rect 495 -1105 545 -1090
rect 575 -555 625 -535
rect 575 -1090 590 -555
rect 610 -1090 625 -555
rect 575 -1105 625 -1090
rect 765 -555 815 -535
rect 765 -1090 780 -555
rect 800 -1090 815 -555
rect 765 -1105 815 -1090
rect 845 -555 895 -535
rect 845 -1090 860 -555
rect 880 -1090 895 -555
rect 845 -1105 895 -1090
rect 1035 -555 1085 -535
rect 1035 -1090 1050 -555
rect 1070 -1090 1085 -555
rect 1035 -1105 1085 -1090
rect 1115 -555 1165 -535
rect 1115 -1090 1130 -555
rect 1150 -1090 1165 -555
rect 1115 -1105 1165 -1090
rect 1305 -555 1355 -535
rect 1305 -1090 1320 -555
rect 1340 -1090 1355 -555
rect 1305 -1105 1355 -1090
rect 1385 -555 1435 -535
rect 1385 -1090 1400 -555
rect 1420 -1090 1435 -555
rect 1385 -1105 1435 -1090
rect 1575 -555 1625 -535
rect 1575 -1090 1590 -555
rect 1610 -1090 1625 -555
rect 1575 -1105 1625 -1090
rect 1655 -555 1705 -535
rect 1655 -1090 1670 -555
rect 1690 -1090 1705 -555
rect 1655 -1105 1705 -1090
rect 1845 -555 1895 -535
rect 1845 -1090 1860 -555
rect 1880 -1090 1895 -555
rect 1845 -1105 1895 -1090
rect 1925 -555 1975 -535
rect 1925 -1090 1940 -555
rect 1960 -1090 1975 -555
rect 1925 -1105 1975 -1090
rect 2115 -555 2165 -535
rect 2115 -1090 2130 -555
rect 2150 -1090 2165 -555
rect 2115 -1105 2165 -1090
rect 2305 -555 2355 -535
rect 2305 -1090 2320 -555
rect 2340 -1090 2355 -555
rect 2305 -1105 2355 -1090
rect 70 -1190 115 -1170
rect 70 -1725 80 -1190
rect 100 -1725 115 -1190
rect 70 -1740 115 -1725
rect 255 -1190 305 -1170
rect 255 -1725 270 -1190
rect 290 -1725 305 -1190
rect 255 -1740 305 -1725
rect 445 -1190 495 -1170
rect 445 -1725 460 -1190
rect 480 -1725 495 -1190
rect 445 -1740 495 -1725
rect 525 -1190 575 -1170
rect 525 -1725 540 -1190
rect 560 -1725 575 -1190
rect 525 -1740 575 -1725
rect 715 -1190 765 -1170
rect 715 -1725 730 -1190
rect 750 -1725 765 -1190
rect 715 -1740 765 -1725
rect 795 -1190 845 -1170
rect 795 -1725 810 -1190
rect 830 -1725 845 -1190
rect 795 -1740 845 -1725
rect 985 -1190 1035 -1170
rect 985 -1725 1000 -1190
rect 1020 -1725 1035 -1190
rect 985 -1740 1035 -1725
rect 1065 -1190 1115 -1170
rect 1065 -1725 1080 -1190
rect 1100 -1725 1115 -1190
rect 1065 -1740 1115 -1725
rect 1255 -1190 1305 -1170
rect 1255 -1725 1270 -1190
rect 1290 -1725 1305 -1190
rect 1255 -1740 1305 -1725
rect 1335 -1190 1385 -1170
rect 1335 -1725 1350 -1190
rect 1370 -1725 1385 -1190
rect 1335 -1740 1385 -1725
rect 1525 -1190 1575 -1170
rect 1525 -1725 1540 -1190
rect 1560 -1725 1575 -1190
rect 1525 -1740 1575 -1725
rect 1605 -1190 1655 -1170
rect 1605 -1725 1620 -1190
rect 1640 -1725 1655 -1190
rect 1605 -1740 1655 -1725
rect 1795 -1190 1845 -1170
rect 1795 -1725 1810 -1190
rect 1830 -1725 1845 -1190
rect 1795 -1740 1845 -1725
rect 1875 -1190 1925 -1170
rect 1875 -1725 1890 -1190
rect 1910 -1725 1925 -1190
rect 1875 -1740 1925 -1725
rect 2065 -1190 2115 -1170
rect 2065 -1725 2080 -1190
rect 2100 -1725 2115 -1190
rect 2065 -1740 2115 -1725
rect 2255 -1190 2305 -1170
rect 2255 -1725 2270 -1190
rect 2290 -1725 2305 -1190
rect 2255 -1740 2305 -1725
<< ndiffc >>
rect -60 -420 -40 115
rect 130 -420 150 115
rect 320 -420 340 115
rect 510 -420 530 115
rect 590 -420 610 115
rect 780 -420 800 115
rect 860 -420 880 115
rect 1050 -420 1070 115
rect 1130 -420 1150 115
rect 1320 -420 1340 115
rect 1400 -420 1420 115
rect 1590 -420 1610 115
rect 1670 -420 1690 115
rect 1860 -420 1880 115
rect 2050 -420 2070 115
rect 130 -1090 150 -555
rect 320 -1090 340 -555
rect 510 -1090 530 -555
rect 590 -1090 610 -555
rect 780 -1090 800 -555
rect 860 -1090 880 -555
rect 1050 -1090 1070 -555
rect 1130 -1090 1150 -555
rect 1320 -1090 1340 -555
rect 1400 -1090 1420 -555
rect 1590 -1090 1610 -555
rect 1670 -1090 1690 -555
rect 1860 -1090 1880 -555
rect 1940 -1090 1960 -555
rect 2130 -1090 2150 -555
rect 2320 -1090 2340 -555
rect 80 -1725 100 -1190
rect 270 -1725 290 -1190
rect 460 -1725 480 -1190
rect 540 -1725 560 -1190
rect 730 -1725 750 -1190
rect 810 -1725 830 -1190
rect 1000 -1725 1020 -1190
rect 1080 -1725 1100 -1190
rect 1270 -1725 1290 -1190
rect 1350 -1725 1370 -1190
rect 1540 -1725 1560 -1190
rect 1620 -1725 1640 -1190
rect 1810 -1725 1830 -1190
rect 1890 -1725 1910 -1190
rect 2080 -1725 2100 -1190
rect 2270 -1725 2290 -1190
<< psubdiff >>
rect 2085 115 2135 135
rect 2085 -420 2100 115
rect 2120 -420 2135 115
rect 2085 -435 2135 -420
rect 70 -555 120 -535
rect 70 -1090 85 -555
rect 105 -1090 120 -555
rect 70 -1105 120 -1090
rect 20 -1190 70 -1170
rect 20 -1725 35 -1190
rect 55 -1725 70 -1190
rect 20 -1740 70 -1725
rect 2305 -1190 2355 -1170
rect 2305 -1725 2320 -1190
rect 2340 -1725 2355 -1190
rect 2305 -1740 2355 -1725
<< psubdiffcont >>
rect 2100 -420 2120 115
rect 85 -1090 105 -555
rect 35 -1725 55 -1190
rect 2320 -1725 2340 -1190
<< poly >>
rect -25 135 115 150
rect 165 135 305 150
rect 355 135 495 150
rect 625 135 765 150
rect 895 135 1035 150
rect 1165 135 1305 150
rect 1435 135 1575 150
rect 1705 135 1845 150
rect 1895 135 2035 150
rect -25 -450 115 -435
rect 165 -445 305 -435
rect 355 -445 495 -435
rect 625 -445 765 -435
rect 895 -445 1035 -435
rect 1165 -445 1305 -435
rect 1435 -445 1575 -435
rect 1705 -445 1845 -435
rect -25 -455 15 -450
rect -25 -475 -15 -455
rect 5 -475 15 -455
rect 165 -460 1845 -445
rect 1895 -450 2035 -435
rect 1995 -455 2035 -450
rect -25 -485 15 -475
rect 165 -495 205 -485
rect 165 -515 175 -495
rect 195 -515 205 -495
rect 165 -520 205 -515
rect 355 -510 445 -460
rect 540 -490 580 -460
rect 540 -510 550 -490
rect 570 -510 580 -490
rect 625 -510 715 -460
rect 810 -490 850 -460
rect 810 -510 820 -490
rect 840 -510 850 -490
rect 895 -510 985 -460
rect 1080 -490 1120 -460
rect 1080 -510 1090 -490
rect 1110 -510 1120 -490
rect 1165 -510 1255 -460
rect 1350 -490 1390 -460
rect 1350 -510 1360 -490
rect 1380 -510 1390 -490
rect 1435 -510 1525 -460
rect 1620 -490 1660 -460
rect 1620 -510 1630 -490
rect 1650 -510 1660 -490
rect 1705 -510 1795 -460
rect 1995 -475 2005 -455
rect 2025 -475 2035 -455
rect 1995 -485 2035 -475
rect 165 -535 305 -520
rect 355 -525 2115 -510
rect 355 -535 495 -525
rect 625 -535 765 -525
rect 895 -535 1035 -525
rect 1165 -535 1305 -525
rect 1435 -535 1575 -525
rect 1705 -535 1845 -525
rect 1975 -535 2115 -525
rect 2165 -535 2305 -520
rect 165 -1120 305 -1105
rect 355 -1115 495 -1105
rect 625 -1115 765 -1105
rect 895 -1115 1035 -1105
rect 1165 -1115 1305 -1105
rect 1435 -1115 1575 -1105
rect 1705 -1115 1845 -1105
rect 1975 -1115 2115 -1105
rect 115 -1130 255 -1120
rect 115 -1150 125 -1130
rect 145 -1150 255 -1130
rect 355 -1130 2115 -1115
rect 2165 -1120 2305 -1105
rect 2165 -1130 2255 -1120
rect 355 -1145 2065 -1130
rect 115 -1170 255 -1150
rect 305 -1160 2065 -1145
rect 2165 -1150 2225 -1130
rect 2245 -1150 2255 -1130
rect 2165 -1155 2255 -1150
rect 305 -1170 445 -1160
rect 575 -1170 715 -1160
rect 845 -1170 985 -1160
rect 1115 -1170 1255 -1160
rect 1385 -1170 1525 -1160
rect 1655 -1170 1795 -1160
rect 1925 -1170 2065 -1160
rect 2115 -1170 2255 -1155
rect 115 -1755 255 -1740
rect 305 -1755 445 -1740
rect 575 -1755 715 -1740
rect 845 -1755 985 -1740
rect 1115 -1755 1255 -1740
rect 1385 -1755 1525 -1740
rect 1655 -1755 1795 -1740
rect 1925 -1755 2065 -1740
rect 2115 -1755 2255 -1740
<< polycont >>
rect -15 -475 5 -455
rect 175 -515 195 -495
rect 550 -510 570 -490
rect 820 -510 840 -490
rect 1090 -510 1110 -490
rect 1360 -510 1380 -490
rect 1630 -510 1650 -490
rect 2005 -475 2025 -455
rect 125 -1150 145 -1130
rect 2225 -1150 2245 -1130
<< locali >>
rect -70 115 -30 130
rect -70 -420 -60 115
rect -40 -420 -30 115
rect -70 -430 -30 -420
rect 120 115 160 130
rect 120 -420 130 115
rect 150 -420 160 115
rect 120 -430 160 -420
rect 310 115 350 130
rect 310 -420 320 115
rect 340 -420 350 115
rect 310 -430 350 -420
rect -50 -445 -30 -430
rect -50 -455 15 -445
rect -50 -465 -15 -455
rect -25 -475 -15 -465
rect 5 -475 15 -455
rect -25 -485 15 -475
rect 165 -495 205 -485
rect 165 -505 175 -495
rect 140 -515 175 -505
rect 195 -515 205 -495
rect 140 -525 205 -515
rect 140 -540 160 -525
rect 330 -540 350 -430
rect 500 115 540 130
rect 500 -420 510 115
rect 530 -420 540 115
rect 500 -430 540 -420
rect 580 115 620 130
rect 580 -420 590 115
rect 610 -420 620 115
rect 580 -430 620 -420
rect 500 -460 520 -430
rect 75 -555 160 -540
rect 75 -1090 85 -555
rect 105 -1090 130 -555
rect 150 -1090 160 -555
rect 75 -1100 160 -1090
rect 310 -555 350 -540
rect 310 -1090 320 -555
rect 340 -1090 350 -555
rect 310 -1100 350 -1090
rect 415 -480 520 -460
rect 310 -1120 330 -1100
rect 115 -1130 155 -1120
rect 115 -1140 125 -1130
rect 90 -1150 125 -1140
rect 145 -1150 155 -1130
rect 90 -1160 155 -1150
rect 280 -1140 330 -1120
rect 415 -1120 435 -480
rect 540 -490 580 -480
rect 540 -500 550 -490
rect 520 -510 550 -500
rect 570 -510 580 -490
rect 520 -520 580 -510
rect 520 -540 540 -520
rect 600 -540 620 -430
rect 770 115 810 130
rect 770 -420 780 115
rect 800 -420 810 115
rect 770 -430 810 -420
rect 850 115 890 130
rect 850 -420 860 115
rect 880 -420 890 115
rect 850 -430 890 -420
rect 770 -460 790 -430
rect 500 -555 540 -540
rect 500 -1090 510 -555
rect 530 -1090 540 -555
rect 500 -1100 540 -1090
rect 580 -555 620 -540
rect 580 -1090 590 -555
rect 610 -1090 620 -555
rect 580 -1100 620 -1090
rect 685 -480 790 -460
rect 580 -1120 600 -1100
rect 415 -1140 470 -1120
rect 90 -1175 110 -1160
rect 280 -1175 300 -1140
rect 25 -1190 110 -1175
rect 25 -1725 35 -1190
rect 55 -1725 80 -1190
rect 100 -1725 110 -1190
rect 25 -1735 110 -1725
rect 260 -1190 300 -1175
rect 260 -1725 270 -1190
rect 290 -1725 300 -1190
rect 260 -1735 300 -1725
rect 450 -1175 470 -1140
rect 550 -1140 600 -1120
rect 685 -1120 705 -480
rect 810 -490 850 -480
rect 810 -500 820 -490
rect 790 -510 820 -500
rect 840 -510 850 -490
rect 790 -520 850 -510
rect 790 -540 810 -520
rect 870 -540 890 -430
rect 1040 115 1080 130
rect 1040 -420 1050 115
rect 1070 -420 1080 115
rect 1040 -430 1080 -420
rect 1120 115 1160 130
rect 1120 -420 1130 115
rect 1150 -420 1160 115
rect 1120 -430 1160 -420
rect 1040 -460 1060 -430
rect 770 -555 810 -540
rect 770 -1090 780 -555
rect 800 -1090 810 -555
rect 770 -1100 810 -1090
rect 850 -555 890 -540
rect 850 -1090 860 -555
rect 880 -1090 890 -555
rect 850 -1100 890 -1090
rect 955 -480 1060 -460
rect 850 -1120 870 -1100
rect 685 -1140 740 -1120
rect 550 -1175 570 -1140
rect 450 -1190 570 -1175
rect 450 -1725 460 -1190
rect 480 -1725 540 -1190
rect 560 -1725 570 -1190
rect 450 -1735 570 -1725
rect 720 -1175 740 -1140
rect 820 -1140 870 -1120
rect 955 -1120 975 -480
rect 1080 -490 1120 -480
rect 1080 -500 1090 -490
rect 1060 -510 1090 -500
rect 1110 -510 1120 -490
rect 1060 -520 1120 -510
rect 1060 -540 1080 -520
rect 1140 -540 1160 -430
rect 1310 115 1350 130
rect 1310 -420 1320 115
rect 1340 -420 1350 115
rect 1310 -430 1350 -420
rect 1390 115 1430 130
rect 1390 -420 1400 115
rect 1420 -420 1430 115
rect 1390 -430 1430 -420
rect 1310 -460 1330 -430
rect 1040 -555 1080 -540
rect 1040 -1090 1050 -555
rect 1070 -1090 1080 -555
rect 1040 -1100 1080 -1090
rect 1120 -555 1160 -540
rect 1120 -1090 1130 -555
rect 1150 -1090 1160 -555
rect 1120 -1100 1160 -1090
rect 1225 -480 1330 -460
rect 1120 -1120 1140 -1100
rect 955 -1140 1010 -1120
rect 820 -1175 840 -1140
rect 720 -1190 840 -1175
rect 720 -1725 730 -1190
rect 750 -1725 810 -1190
rect 830 -1725 840 -1190
rect 720 -1735 840 -1725
rect 990 -1175 1010 -1140
rect 1090 -1140 1140 -1120
rect 1225 -1120 1245 -480
rect 1350 -490 1390 -480
rect 1350 -500 1360 -490
rect 1330 -510 1360 -500
rect 1380 -510 1390 -490
rect 1330 -520 1390 -510
rect 1330 -540 1350 -520
rect 1410 -540 1430 -430
rect 1580 115 1620 130
rect 1580 -420 1590 115
rect 1610 -420 1620 115
rect 1580 -430 1620 -420
rect 1660 115 1700 130
rect 1660 -420 1670 115
rect 1690 -420 1700 115
rect 1660 -430 1700 -420
rect 1580 -460 1600 -430
rect 1310 -555 1350 -540
rect 1310 -1090 1320 -555
rect 1340 -1090 1350 -555
rect 1310 -1100 1350 -1090
rect 1390 -555 1430 -540
rect 1390 -1090 1400 -555
rect 1420 -1090 1430 -555
rect 1390 -1100 1430 -1090
rect 1495 -480 1600 -460
rect 1390 -1120 1410 -1100
rect 1225 -1140 1280 -1120
rect 1090 -1175 1110 -1140
rect 990 -1190 1110 -1175
rect 990 -1725 1000 -1190
rect 1020 -1725 1080 -1190
rect 1100 -1725 1110 -1190
rect 990 -1735 1110 -1725
rect 1260 -1175 1280 -1140
rect 1360 -1140 1410 -1120
rect 1495 -1120 1515 -480
rect 1620 -490 1660 -480
rect 1620 -500 1630 -490
rect 1600 -510 1630 -500
rect 1650 -510 1660 -490
rect 1600 -520 1660 -510
rect 1600 -540 1620 -520
rect 1680 -540 1700 -430
rect 1850 115 1890 130
rect 1850 -420 1860 115
rect 1880 -420 1890 115
rect 1850 -430 1890 -420
rect 2040 115 2130 130
rect 2040 -420 2050 115
rect 2070 -420 2100 115
rect 2120 -420 2130 115
rect 2040 -430 2130 -420
rect 1850 -460 1870 -430
rect 2040 -445 2060 -430
rect 1580 -555 1620 -540
rect 1580 -1090 1590 -555
rect 1610 -1090 1620 -555
rect 1580 -1100 1620 -1090
rect 1660 -555 1700 -540
rect 1660 -1090 1670 -555
rect 1690 -1090 1700 -555
rect 1660 -1100 1700 -1090
rect 1765 -480 1870 -460
rect 1995 -455 2060 -445
rect 1995 -475 2005 -455
rect 2025 -465 2060 -455
rect 2025 -475 2035 -465
rect 1660 -1120 1680 -1100
rect 1495 -1140 1550 -1120
rect 1360 -1175 1380 -1140
rect 1260 -1190 1380 -1175
rect 1260 -1725 1270 -1190
rect 1290 -1725 1350 -1190
rect 1370 -1725 1380 -1190
rect 1260 -1735 1380 -1725
rect 1530 -1175 1550 -1140
rect 1630 -1140 1680 -1120
rect 1765 -1120 1785 -480
rect 1995 -485 2035 -475
rect 2140 -485 2355 -465
rect 2140 -540 2160 -485
rect 1850 -555 1890 -540
rect 1850 -1090 1860 -555
rect 1880 -1090 1890 -555
rect 1850 -1100 1890 -1090
rect 1930 -555 1970 -540
rect 1930 -1090 1940 -555
rect 1960 -1090 1970 -555
rect 1930 -1100 1970 -1090
rect 2120 -555 2160 -540
rect 2120 -1090 2130 -555
rect 2150 -1090 2160 -555
rect 2120 -1100 2160 -1090
rect 2310 -555 2350 -540
rect 2310 -1090 2320 -555
rect 2340 -1090 2350 -555
rect 2310 -1100 2350 -1090
rect 1930 -1120 1950 -1100
rect 2120 -1120 2140 -1100
rect 1765 -1140 1820 -1120
rect 1630 -1175 1650 -1140
rect 1530 -1190 1650 -1175
rect 1530 -1725 1540 -1190
rect 1560 -1725 1620 -1190
rect 1640 -1725 1650 -1190
rect 1530 -1735 1650 -1725
rect 1800 -1175 1820 -1140
rect 1900 -1140 1950 -1120
rect 2090 -1140 2140 -1120
rect 2215 -1130 2255 -1120
rect 1900 -1175 1920 -1140
rect 2090 -1175 2110 -1140
rect 2215 -1150 2225 -1130
rect 2245 -1140 2255 -1130
rect 2245 -1150 2280 -1140
rect 2215 -1160 2280 -1150
rect 1800 -1190 1920 -1175
rect 1800 -1725 1810 -1190
rect 1830 -1725 1890 -1190
rect 1910 -1725 1920 -1190
rect 1800 -1735 1920 -1725
rect 2070 -1190 2110 -1175
rect 2070 -1725 2080 -1190
rect 2100 -1725 2110 -1190
rect 2070 -1735 2110 -1725
rect 2260 -1175 2280 -1160
rect 2260 -1190 2350 -1175
rect 2260 -1725 2270 -1190
rect 2290 -1725 2320 -1190
rect 2340 -1725 2350 -1190
rect 2260 -1735 2350 -1725
rect 280 -1780 300 -1735
rect 550 -1780 570 -1735
rect 820 -1780 840 -1735
rect 1090 -1780 1110 -1735
rect 1360 -1780 1380 -1735
rect 1630 -1780 1650 -1735
rect 1900 -1780 1920 -1735
<< viali >>
rect -60 -420 -40 115
rect 130 -420 150 -370
rect 85 -1090 105 -555
rect 130 -1090 150 -555
rect 510 -605 530 -555
rect 35 -1725 55 -1190
rect 80 -1725 100 -1190
rect 780 -605 800 -555
rect 1050 -605 1070 -555
rect 1320 -605 1340 -555
rect 2050 -420 2070 115
rect 2100 -420 2120 115
rect 1590 -605 1610 -555
rect 1860 -605 1880 -555
rect 2320 -1090 2340 -555
rect 2270 -1725 2290 -1190
rect 2320 -1725 2340 -1190
<< metal1 >>
rect -75 115 2150 130
rect -75 -420 -60 115
rect -40 -315 2050 115
rect -40 -420 -30 -315
rect -75 -430 -30 -420
rect -15 -370 540 -345
rect -15 -420 130 -370
rect 150 -420 540 -370
rect -15 -425 540 -420
rect -15 -535 40 -425
rect -75 -730 40 -535
rect 500 -540 540 -425
rect 580 -420 2050 -315
rect 2070 -420 2100 115
rect 2120 -420 2150 115
rect 580 -430 2150 -420
rect 2040 -540 2150 -430
rect 75 -555 160 -540
rect 75 -1090 85 -555
rect 105 -1090 130 -555
rect 150 -650 160 -555
rect 500 -555 1890 -540
rect 500 -605 510 -555
rect 530 -605 780 -555
rect 800 -605 1050 -555
rect 1070 -605 1320 -555
rect 1340 -605 1590 -555
rect 1610 -605 1860 -555
rect 1880 -605 1890 -555
rect 500 -620 1890 -605
rect 1930 -555 2350 -540
rect 1930 -650 2320 -555
rect 150 -1090 2320 -650
rect 2340 -1090 2350 -555
rect 75 -1175 2350 -1090
rect -75 -1190 2350 -1175
rect -75 -1725 35 -1190
rect 55 -1725 80 -1190
rect 100 -1725 2270 -1190
rect 2290 -1725 2320 -1190
rect 2340 -1725 2350 -1190
rect -75 -1735 2350 -1725
<< labels >>
rlabel metal1 -75 -630 -75 -630 7 VP
rlabel metal1 -75 -1455 -75 -1455 7 VN
rlabel locali 2355 -475 2355 -475 3 Iout
rlabel locali 290 -1780 290 -1780 5 branch0
rlabel locali 560 -1780 560 -1780 5 branch1
rlabel locali 830 -1780 830 -1780 5 branch2
rlabel locali 1100 -1780 1100 -1780 5 branch3
rlabel locali 1370 -1780 1370 -1780 5 branch4
rlabel locali 1640 -1780 1640 -1780 5 branch5
rlabel locali 1910 -1780 1910 -1780 5 branch6
<< end >>
