* SPICE3 file created from biasgen.ext - technology: sky130A


* Top level circuit biasgen

X0 a_50_260# a_50_n170# VP VP sky130_fd_pr__pfet_01v8 ad=3.5e+11p pd=2.4e+06u as=5.25e+12p ps=3.6e+07u w=700000u l=500000u
X1 VN VN a_50_260# VN sky130_fd_pr__nfet_01v8 ad=1.085e+13p pd=6.04e+07u as=7e+11p ps=4.8e+06u w=700000u l=500000u
X2 a_n30_n580# VN VN VN sky130_fd_pr__nfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X3 a_n430_n580# a_n430_n580# VP VP sky130_fd_pr__pfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X4 a_50_n170# VN VN VN sky130_fd_pr__nfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X5 VN a_n30_n580# a_570_n1030# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.05e+12p ps=7.2e+06u w=700000u l=500000u
X6 VP a_n430_n580# a_n430_n580# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X7 a_n1050_n90# VN VN VN sky130_fd_pr__nfet_01v8 ad=5.6e+12p pd=2.44e+07u as=0p ps=0u w=5.6e+06u l=500000u
X8 Rbias a_n1050_n90# a_n1050_n90# VN sky130_fd_pr__nfet_01v8 ad=2.8e+12p pd=1.22e+07u as=0p ps=0u w=5.6e+06u l=500000u
X9 a_50_n170# VP VP VP sky130_fd_pr__pfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X10 a_50_260# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X11 a_570_n1030# a_n30_n580# a_n30_n580# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X12 a_n1050_n90# a_50_260# VP VP sky130_fd_pr__pfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X13 VN Vbn Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5e+11p ps=2.4e+06u w=700000u l=500000u
X14 VN VN a_50_n170# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X15 VP a_50_260# Vbn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.5e+11p ps=2.4e+06u w=700000u l=500000u
X16 Vc Vc a_570_n1030# VN sky130_fd_pr__nfet_01v8 ad=3.5e+11p pd=2.4e+06u as=0p ps=0u w=700000u l=500000u
X17 Vc a_50_260# VP VP sky130_fd_pr__pfet_01v8 ad=3.5e+11p pd=2.4e+06u as=0p ps=0u w=700000u l=500000u
X18 VN Rbias a_n430_n580# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5e+11p ps=2.4e+06u w=700000u l=500000u
X19 VN VN a_n1050_n90# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.6e+06u l=500000u
X20 a_570_n1030# Vc Vc VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X21 VN Vbn a_50_260# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X22 a_n30_n580# a_n430_n580# VP VP sky130_fd_pr__pfet_01v8 ad=3.5e+11p pd=2.4e+06u as=0p ps=0u w=700000u l=500000u
X23 a_n430_n580# Rbias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X24 VP a_50_260# a_n1050_n90# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X25 a_50_n170# a_50_n170# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X26 VP a_50_n170# a_50_260# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X27 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X28 a_50_n170# a_n1050_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X29 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X30 VP a_n430_n580# a_n30_n580# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X31 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X32 VP a_50_n170# a_50_n170# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X33 VP VP a_n1050_n90# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X34 a_50_260# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X35 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X36 a_570_n1030# a_n30_n580# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X37 VP a_50_260# Vc VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X38 VN a_n1050_n90# a_50_n170# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X39 a_n1050_n90# a_n1050_n90# Rbias VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.6e+06u l=500000u
X40 Vbn Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X41 a_n30_n580# a_n30_n580# a_570_n1030# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X42 Vbn a_50_260# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X43 VP VP a_50_n170# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X44 VP VP a_n430_n580# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X45 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X46 a_n430_n580# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X47 VN VN a_n30_n580# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X48 a_n1050_n90# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X49 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
.end

