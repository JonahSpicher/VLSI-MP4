magic
tech sky130A
timestamp 1618368219
<< nwell >>
rect 5 285 745 570
rect -385 -310 755 -195
<< nmos >>
rect -575 -45 -525 515
rect -475 -45 -425 515
rect -375 -45 -325 515
rect -275 -45 -225 515
rect -25 130 25 200
rect 75 130 125 200
rect 175 130 225 200
rect 275 130 325 200
rect 375 130 425 200
rect 475 130 525 200
rect -25 -85 25 -15
rect 75 -85 125 -15
rect 175 -85 225 -15
rect 275 -85 325 -15
rect 375 -85 425 -15
rect 475 -85 525 -15
rect 575 -85 625 -15
rect 675 -85 725 -15
rect -265 -515 -215 -445
rect -165 -515 -115 -445
rect -65 -515 -15 -445
rect 35 -515 85 -445
rect 135 -515 185 -445
rect 235 -515 285 -445
rect 335 -515 385 -445
rect 435 -515 485 -445
rect 535 -515 585 -445
rect 635 -515 685 -445
<< pmos >>
rect 125 480 175 550
rect 225 480 275 550
rect 325 480 375 550
rect 425 480 475 550
rect 525 480 575 550
rect 625 480 675 550
rect 125 305 175 375
rect 225 305 275 375
rect 325 305 375 375
rect 425 305 475 375
rect 525 305 575 375
rect 625 305 675 375
rect -265 -290 -215 -220
rect -165 -290 -115 -220
rect -65 -290 -15 -220
rect 35 -290 85 -220
rect 135 -290 185 -220
rect 235 -290 285 -220
rect 335 -290 385 -220
rect 435 -290 485 -220
rect 535 -290 585 -220
rect 635 -290 685 -220
<< ndiff >>
rect -625 500 -575 515
rect -625 -30 -610 500
rect -590 -30 -575 500
rect -625 -45 -575 -30
rect -525 500 -475 515
rect -525 -30 -510 500
rect -490 -30 -475 500
rect -525 -45 -475 -30
rect -425 500 -375 515
rect -425 -30 -410 500
rect -390 -30 -375 500
rect -425 -45 -375 -30
rect -325 500 -275 515
rect -325 -30 -310 500
rect -290 -30 -275 500
rect -325 -45 -275 -30
rect -225 500 -175 515
rect -225 -30 -210 500
rect -190 -30 -175 500
rect -75 185 -25 200
rect -75 145 -60 185
rect -40 145 -25 185
rect -75 130 -25 145
rect 25 185 75 200
rect 25 145 40 185
rect 60 145 75 185
rect 25 130 75 145
rect 125 185 175 200
rect 125 145 140 185
rect 160 145 175 185
rect 125 130 175 145
rect 225 185 275 200
rect 225 145 240 185
rect 260 145 275 185
rect 225 130 275 145
rect 325 185 375 200
rect 325 145 340 185
rect 360 145 375 185
rect 325 130 375 145
rect 425 185 475 200
rect 425 145 440 185
rect 460 145 475 185
rect 425 130 475 145
rect 525 185 575 200
rect 525 145 540 185
rect 560 145 575 185
rect 525 130 575 145
rect -225 -45 -175 -30
rect -75 -30 -25 -15
rect -75 -70 -60 -30
rect -40 -70 -25 -30
rect -75 -85 -25 -70
rect 25 -30 75 -15
rect 25 -70 40 -30
rect 60 -70 75 -30
rect 25 -85 75 -70
rect 125 -30 175 -15
rect 125 -70 140 -30
rect 160 -70 175 -30
rect 125 -85 175 -70
rect 225 -30 275 -15
rect 225 -70 240 -30
rect 260 -70 275 -30
rect 225 -85 275 -70
rect 325 -30 375 -15
rect 325 -70 340 -30
rect 360 -70 375 -30
rect 325 -85 375 -70
rect 425 -30 475 -15
rect 425 -70 440 -30
rect 460 -70 475 -30
rect 425 -85 475 -70
rect 525 -30 575 -15
rect 525 -70 540 -30
rect 560 -70 575 -30
rect 525 -85 575 -70
rect 625 -30 675 -15
rect 625 -70 640 -30
rect 660 -70 675 -30
rect 625 -85 675 -70
rect 725 -30 775 -15
rect 725 -70 740 -30
rect 760 -70 775 -30
rect 725 -85 775 -70
rect -315 -460 -265 -445
rect -315 -500 -300 -460
rect -280 -500 -265 -460
rect -315 -515 -265 -500
rect -215 -460 -165 -445
rect -215 -500 -200 -460
rect -180 -500 -165 -460
rect -215 -515 -165 -500
rect -115 -460 -65 -445
rect -115 -500 -100 -460
rect -80 -500 -65 -460
rect -115 -515 -65 -500
rect -15 -460 35 -445
rect -15 -500 0 -460
rect 20 -500 35 -460
rect -15 -515 35 -500
rect 85 -460 135 -445
rect 85 -500 100 -460
rect 120 -500 135 -460
rect 85 -515 135 -500
rect 185 -460 235 -445
rect 185 -500 200 -460
rect 220 -500 235 -460
rect 185 -515 235 -500
rect 285 -460 335 -445
rect 285 -500 300 -460
rect 320 -500 335 -460
rect 285 -515 335 -500
rect 385 -460 435 -445
rect 385 -500 400 -460
rect 420 -500 435 -460
rect 385 -515 435 -500
rect 485 -460 535 -445
rect 485 -500 500 -460
rect 520 -500 535 -460
rect 485 -515 535 -500
rect 585 -460 635 -445
rect 585 -500 600 -460
rect 620 -500 635 -460
rect 585 -515 635 -500
rect 685 -460 735 -445
rect 685 -500 700 -460
rect 720 -500 735 -460
rect 685 -515 735 -500
<< pdiff >>
rect 75 535 125 550
rect 75 495 90 535
rect 110 495 125 535
rect 75 480 125 495
rect 175 535 225 550
rect 175 495 190 535
rect 210 495 225 535
rect 175 480 225 495
rect 275 535 325 550
rect 275 495 290 535
rect 310 495 325 535
rect 275 480 325 495
rect 375 535 425 550
rect 375 495 390 535
rect 410 495 425 535
rect 375 480 425 495
rect 475 535 525 550
rect 475 495 490 535
rect 510 495 525 535
rect 475 480 525 495
rect 575 535 625 550
rect 575 495 590 535
rect 610 495 625 535
rect 575 480 625 495
rect 675 535 725 550
rect 675 495 690 535
rect 710 495 725 535
rect 675 480 725 495
rect 75 360 125 375
rect 75 320 90 360
rect 110 320 125 360
rect 75 305 125 320
rect 175 360 225 375
rect 175 320 190 360
rect 210 320 225 360
rect 175 305 225 320
rect 275 360 325 375
rect 275 320 290 360
rect 310 320 325 360
rect 275 305 325 320
rect 375 360 425 375
rect 375 320 390 360
rect 410 320 425 360
rect 375 305 425 320
rect 475 360 525 375
rect 475 320 490 360
rect 510 320 525 360
rect 475 305 525 320
rect 575 360 625 375
rect 575 320 590 360
rect 610 320 625 360
rect 575 305 625 320
rect 675 360 725 375
rect 675 320 690 360
rect 710 320 725 360
rect 675 305 725 320
rect -315 -235 -265 -220
rect -315 -275 -300 -235
rect -280 -275 -265 -235
rect -315 -290 -265 -275
rect -215 -235 -165 -220
rect -215 -275 -200 -235
rect -180 -275 -165 -235
rect -215 -290 -165 -275
rect -115 -235 -65 -220
rect -115 -275 -100 -235
rect -80 -275 -65 -235
rect -115 -290 -65 -275
rect -15 -235 35 -220
rect -15 -275 0 -235
rect 20 -275 35 -235
rect -15 -290 35 -275
rect 85 -235 135 -220
rect 85 -275 100 -235
rect 120 -275 135 -235
rect 85 -290 135 -275
rect 185 -235 235 -220
rect 185 -275 200 -235
rect 220 -275 235 -235
rect 185 -290 235 -275
rect 285 -235 335 -220
rect 285 -275 300 -235
rect 320 -275 335 -235
rect 285 -290 335 -275
rect 385 -235 435 -220
rect 385 -275 400 -235
rect 420 -275 435 -235
rect 385 -290 435 -275
rect 485 -235 535 -220
rect 485 -275 500 -235
rect 520 -275 535 -235
rect 485 -290 535 -275
rect 585 -235 635 -220
rect 585 -275 600 -235
rect 620 -275 635 -235
rect 585 -290 635 -275
rect 685 -235 735 -220
rect 685 -275 700 -235
rect 720 -275 735 -235
rect 685 -290 735 -275
<< ndiffc >>
rect -610 -30 -590 500
rect -510 -30 -490 500
rect -410 -30 -390 500
rect -310 -30 -290 500
rect -210 -30 -190 500
rect -60 145 -40 185
rect 40 145 60 185
rect 140 145 160 185
rect 240 145 260 185
rect 340 145 360 185
rect 440 145 460 185
rect 540 145 560 185
rect -60 -70 -40 -30
rect 40 -70 60 -30
rect 140 -70 160 -30
rect 240 -70 260 -30
rect 340 -70 360 -30
rect 440 -70 460 -30
rect 540 -70 560 -30
rect 640 -70 660 -30
rect 740 -70 760 -30
rect -300 -500 -280 -460
rect -200 -500 -180 -460
rect -100 -500 -80 -460
rect 0 -500 20 -460
rect 100 -500 120 -460
rect 200 -500 220 -460
rect 300 -500 320 -460
rect 400 -500 420 -460
rect 500 -500 520 -460
rect 600 -500 620 -460
rect 700 -500 720 -460
<< pdiffc >>
rect 90 495 110 535
rect 190 495 210 535
rect 290 495 310 535
rect 390 495 410 535
rect 490 495 510 535
rect 590 495 610 535
rect 690 495 710 535
rect 90 320 110 360
rect 190 320 210 360
rect 290 320 310 360
rect 390 320 410 360
rect 490 320 510 360
rect 590 320 610 360
rect 690 320 710 360
rect -300 -275 -280 -235
rect -200 -275 -180 -235
rect -100 -275 -80 -235
rect 0 -275 20 -235
rect 100 -275 120 -235
rect 200 -275 220 -235
rect 300 -275 320 -235
rect 400 -275 420 -235
rect 500 -275 520 -235
rect 600 -275 620 -235
rect 700 -275 720 -235
<< psubdiff >>
rect -125 185 -75 200
rect -125 145 -110 185
rect -90 145 -75 185
rect -125 130 -75 145
rect -365 -460 -315 -445
rect -365 -500 -350 -460
rect -330 -500 -315 -460
rect -365 -515 -315 -500
<< nsubdiff >>
rect 25 535 75 550
rect 25 495 40 535
rect 60 495 75 535
rect 25 480 75 495
rect 25 360 75 375
rect 25 320 40 360
rect 60 320 75 360
rect 25 305 75 320
rect -365 -235 -315 -220
rect -365 -275 -350 -235
rect -330 -275 -315 -235
rect -365 -290 -315 -275
<< psubdiffcont >>
rect -110 145 -90 185
rect -350 -500 -330 -460
<< nsubdiffcont >>
rect 40 495 60 535
rect 40 320 60 360
rect -350 -275 -330 -235
<< poly >>
rect 635 595 675 605
rect 635 575 645 595
rect 665 575 675 595
rect -575 555 -535 565
rect -575 535 -565 555
rect -545 535 -535 555
rect -365 555 -325 565
rect -365 540 -355 555
rect -575 530 -535 535
rect -475 535 -355 540
rect -335 535 -325 555
rect -575 515 -525 530
rect -475 525 -325 535
rect -265 555 -225 565
rect -265 535 -255 555
rect -235 535 -225 555
rect 125 550 175 565
rect 225 560 575 575
rect 635 565 675 575
rect 225 550 275 560
rect 325 550 375 560
rect 425 550 475 560
rect 525 550 575 560
rect 625 550 675 565
rect -265 530 -225 535
rect -475 515 -425 525
rect -375 515 -325 525
rect -275 515 -225 530
rect 125 465 175 480
rect 225 465 275 480
rect 325 465 375 480
rect 425 465 475 480
rect 525 465 575 480
rect 625 465 675 480
rect 125 455 165 465
rect 125 435 135 455
rect 155 435 165 455
rect 325 455 365 465
rect 325 435 335 455
rect 355 435 365 455
rect 50 420 90 430
rect 125 425 165 435
rect 225 425 265 435
rect 325 425 365 435
rect 50 400 60 420
rect 80 400 90 420
rect 225 415 235 425
rect 220 405 235 415
rect 255 405 265 425
rect 220 400 265 405
rect 50 385 175 400
rect 220 395 575 400
rect 125 375 175 385
rect 225 385 575 395
rect 225 375 275 385
rect 325 375 375 385
rect 425 375 475 385
rect 525 375 575 385
rect 625 375 675 390
rect 125 290 175 305
rect 225 290 275 305
rect 325 290 375 305
rect 425 290 475 305
rect 525 290 575 305
rect 625 290 675 305
rect 560 265 575 290
rect 660 265 675 290
rect 560 255 610 265
rect 560 250 580 255
rect -25 240 15 250
rect -25 220 -15 240
rect 5 220 15 240
rect 230 240 270 250
rect 230 225 240 240
rect -25 215 15 220
rect 75 220 240 225
rect 260 225 270 240
rect 485 240 525 250
rect 260 220 425 225
rect -25 200 25 215
rect 75 210 425 220
rect 485 220 495 240
rect 515 220 525 240
rect 570 235 580 250
rect 600 235 610 255
rect 570 225 610 235
rect 635 255 675 265
rect 635 235 645 255
rect 665 235 675 255
rect 635 225 675 235
rect 485 215 525 220
rect 75 200 125 210
rect 175 200 225 210
rect 275 200 325 210
rect 375 200 425 210
rect 475 200 525 215
rect -25 115 25 130
rect 75 115 125 130
rect 175 115 225 130
rect 275 115 325 130
rect 375 115 425 130
rect 475 115 525 130
rect 760 105 800 115
rect 760 85 770 105
rect 790 85 800 105
rect 760 75 800 85
rect -135 60 90 75
rect -135 35 -120 60
rect -155 25 -115 35
rect -155 5 -145 25
rect -125 5 -115 25
rect -155 -5 -115 5
rect -25 25 15 35
rect -25 5 -15 25
rect 5 5 15 25
rect -25 0 15 5
rect 75 15 90 60
rect 330 30 370 40
rect 330 15 340 30
rect 75 0 225 15
rect -25 -15 25 0
rect 75 -15 125 0
rect 175 -15 225 0
rect 275 10 340 15
rect 360 15 370 30
rect 685 30 725 40
rect 360 10 425 15
rect 275 0 425 10
rect 275 -15 325 0
rect 375 -15 425 0
rect 475 0 625 15
rect 685 10 695 30
rect 715 10 725 30
rect 685 5 725 10
rect 475 -15 525 0
rect 575 -15 625 0
rect 675 -15 725 5
rect -575 -60 -525 -45
rect -475 -60 -425 -45
rect -375 -60 -325 -45
rect -275 -60 -225 -45
rect -25 -100 25 -85
rect 75 -100 125 -85
rect 175 -100 225 -85
rect 275 -100 325 -85
rect 375 -100 425 -85
rect 475 -100 525 -85
rect 575 -100 625 -85
rect 675 -100 725 -85
rect 475 -125 490 -100
rect 785 -125 800 75
rect -10 -140 490 -125
rect 570 -140 800 -125
rect -10 -160 0 -140
rect 20 -160 30 -140
rect -265 -175 -225 -165
rect -265 -195 -255 -175
rect -235 -195 -225 -175
rect -265 -205 -225 -195
rect -165 -175 -125 -165
rect -10 -170 30 -160
rect -165 -195 -155 -175
rect -135 -195 -125 -175
rect 145 -175 185 -165
rect 145 -195 155 -175
rect 175 -195 185 -175
rect 290 -175 330 -165
rect 290 -195 300 -175
rect 320 -195 330 -175
rect 570 -195 585 -140
rect -265 -220 -215 -205
rect -165 -210 185 -195
rect -165 -220 -115 -210
rect -65 -220 -15 -210
rect 35 -220 85 -210
rect 135 -220 185 -210
rect 235 -210 385 -195
rect 235 -220 285 -210
rect 335 -220 385 -210
rect 435 -210 585 -195
rect 645 -175 685 -165
rect 645 -195 655 -175
rect 675 -195 685 -175
rect 645 -205 685 -195
rect 435 -220 485 -210
rect 535 -220 585 -210
rect 635 -220 685 -205
rect 745 -185 785 -175
rect 745 -205 755 -185
rect 775 -205 785 -185
rect 745 -215 785 -205
rect -265 -305 -215 -290
rect -165 -305 -115 -290
rect -65 -305 -15 -290
rect 35 -305 85 -290
rect 135 -305 185 -290
rect 235 -305 285 -290
rect 335 -305 385 -290
rect 435 -305 485 -290
rect 535 -305 585 -290
rect 635 -305 685 -290
rect -325 -340 -285 -330
rect -325 -360 -315 -340
rect -295 -355 -285 -340
rect 745 -355 760 -215
rect -295 -360 -150 -355
rect -325 -370 -150 -360
rect -265 -405 -225 -395
rect -265 -425 -255 -405
rect -235 -425 -225 -405
rect -265 -430 -225 -425
rect -165 -420 -150 -370
rect 490 -365 530 -355
rect 490 -380 500 -365
rect 470 -385 500 -380
rect 520 -385 530 -365
rect 470 -395 530 -385
rect 740 -365 780 -355
rect 740 -385 750 -365
rect 770 -385 780 -365
rect 740 -395 780 -385
rect 90 -405 130 -395
rect 90 -420 100 -405
rect -265 -445 -215 -430
rect -165 -435 -15 -420
rect -165 -445 -115 -435
rect -65 -445 -15 -435
rect 35 -425 100 -420
rect 120 -420 130 -405
rect 390 -405 430 -395
rect 390 -420 400 -405
rect 120 -425 185 -420
rect 35 -435 185 -425
rect 335 -425 400 -420
rect 420 -420 430 -405
rect 470 -420 485 -395
rect 420 -425 485 -420
rect 35 -445 85 -435
rect 135 -445 185 -435
rect 235 -445 285 -430
rect 335 -435 485 -425
rect 645 -405 685 -395
rect 645 -425 655 -405
rect 675 -425 685 -405
rect 645 -430 685 -425
rect 335 -445 385 -435
rect 435 -445 485 -435
rect 535 -445 585 -430
rect 635 -445 685 -430
rect -265 -530 -215 -515
rect -165 -530 -115 -515
rect -65 -530 -15 -515
rect 35 -530 85 -515
rect 135 -530 185 -515
rect 235 -530 285 -515
rect 335 -530 385 -515
rect 435 -530 485 -515
rect 535 -530 585 -515
rect 635 -530 685 -515
rect 235 -535 275 -530
rect 235 -555 245 -535
rect 265 -555 275 -535
rect 235 -565 275 -555
rect 545 -535 585 -530
rect 545 -555 555 -535
rect 575 -555 585 -535
rect 545 -565 585 -555
<< polycont >>
rect 645 575 665 595
rect -565 535 -545 555
rect -355 535 -335 555
rect -255 535 -235 555
rect 135 435 155 455
rect 335 435 355 455
rect 60 400 80 420
rect 235 405 255 425
rect -15 220 5 240
rect 240 220 260 240
rect 495 220 515 240
rect 580 235 600 255
rect 645 235 665 255
rect 770 85 790 105
rect -145 5 -125 25
rect -15 5 5 25
rect 340 10 360 30
rect 695 10 715 30
rect 0 -160 20 -140
rect -255 -195 -235 -175
rect -155 -195 -135 -175
rect 155 -195 175 -175
rect 300 -195 320 -175
rect 655 -195 675 -175
rect 755 -205 775 -185
rect -315 -360 -295 -340
rect -255 -425 -235 -405
rect 500 -385 520 -365
rect 750 -385 770 -365
rect 100 -425 120 -405
rect 400 -425 420 -405
rect 655 -425 675 -405
rect 245 -555 265 -535
rect 555 -555 575 -535
<< locali >>
rect -345 585 200 605
rect 635 595 675 605
rect -345 565 -325 585
rect 180 565 600 585
rect 635 575 645 595
rect 665 585 675 595
rect 665 575 700 585
rect 635 565 700 575
rect -575 555 -535 565
rect -575 545 -565 555
rect -600 535 -565 545
rect -545 535 -535 555
rect -365 555 -325 565
rect -365 550 -355 555
rect -600 525 -535 535
rect -500 535 -355 550
rect -335 545 -325 555
rect -265 555 -225 565
rect -335 535 -300 545
rect -500 530 -300 535
rect -600 510 -580 525
rect -500 510 -480 530
rect -365 525 -300 530
rect -265 535 -255 555
rect -235 545 -225 555
rect 180 545 200 565
rect 580 545 600 565
rect 680 545 700 565
rect -235 535 -200 545
rect -265 525 -200 535
rect -320 510 -300 525
rect -220 510 -200 525
rect 30 535 120 545
rect -620 500 -580 510
rect -620 -30 -610 500
rect -590 -30 -580 500
rect -620 -40 -580 -30
rect -520 500 -480 510
rect -520 -30 -510 500
rect -490 -30 -480 500
rect -520 -40 -480 -30
rect -420 500 -380 510
rect -420 -30 -410 500
rect -390 -30 -380 500
rect -420 -40 -380 -30
rect -320 500 -280 510
rect -320 -30 -310 500
rect -290 -30 -280 500
rect -320 -40 -280 -30
rect -220 500 -180 510
rect -220 -30 -210 500
rect -190 -30 -180 500
rect 30 495 40 535
rect 60 495 90 535
rect 110 495 120 535
rect 30 485 120 495
rect 180 535 220 545
rect 180 495 190 535
rect 210 495 220 535
rect 180 485 220 495
rect 280 535 320 545
rect 280 495 290 535
rect 310 495 320 535
rect 280 485 320 495
rect 380 535 420 545
rect 380 495 390 535
rect 410 495 420 535
rect 380 485 420 495
rect 480 535 520 545
rect 480 495 490 535
rect 510 495 520 535
rect 480 485 520 495
rect 580 535 620 545
rect 580 495 590 535
rect 610 495 620 535
rect 580 485 620 495
rect 680 535 720 545
rect 680 495 690 535
rect 710 495 720 535
rect 680 485 720 495
rect 100 465 120 485
rect 400 465 420 485
rect 100 455 165 465
rect 100 445 135 455
rect 125 435 135 445
rect 155 435 165 455
rect 325 455 365 465
rect 325 435 335 455
rect 355 435 365 455
rect 400 455 755 465
rect 400 445 705 455
rect 50 420 90 430
rect 125 425 165 435
rect 225 425 265 435
rect 325 425 365 435
rect 690 435 705 445
rect 740 435 755 455
rect 690 425 755 435
rect 50 400 60 420
rect 80 400 90 420
rect 225 415 235 425
rect 50 370 90 400
rect 200 405 235 415
rect 255 405 265 425
rect 200 395 265 405
rect 335 400 355 425
rect 200 370 220 395
rect 335 380 400 400
rect 380 370 400 380
rect 30 360 120 370
rect 30 320 40 360
rect 60 320 90 360
rect 110 320 120 360
rect 30 310 120 320
rect 180 360 220 370
rect 180 320 190 360
rect 210 320 220 360
rect 180 310 220 320
rect 280 360 320 370
rect 280 320 290 360
rect 310 320 320 360
rect 280 310 320 320
rect 380 360 420 370
rect 380 320 390 360
rect 410 320 420 360
rect 380 310 420 320
rect 480 360 520 370
rect 480 320 490 360
rect 510 320 520 360
rect 480 310 520 320
rect 580 360 620 370
rect 580 320 590 360
rect 610 320 620 360
rect 580 310 620 320
rect 680 360 720 370
rect 680 320 690 360
rect 710 320 720 360
rect 680 310 720 320
rect 180 290 200 310
rect -160 270 200 290
rect 400 275 420 310
rect -160 75 -140 270
rect 230 255 270 265
rect 400 255 450 275
rect 580 265 600 310
rect 680 265 700 310
rect -25 240 15 250
rect -25 230 -15 240
rect -50 220 -15 230
rect 5 220 15 240
rect -50 210 15 220
rect 230 220 240 255
rect 260 220 270 255
rect -50 195 -30 210
rect -120 185 -30 195
rect -120 145 -110 185
rect -90 145 -60 185
rect -40 145 -30 185
rect -120 135 -30 145
rect 30 185 70 195
rect 30 145 40 185
rect 60 145 70 185
rect 30 135 70 145
rect 130 185 170 195
rect 130 145 140 185
rect 160 145 170 185
rect 130 135 170 145
rect 230 185 270 220
rect 430 195 450 255
rect 570 255 610 265
rect 485 240 525 250
rect 485 220 495 240
rect 515 230 525 240
rect 570 235 580 255
rect 600 235 610 255
rect 515 220 550 230
rect 570 225 610 235
rect 635 255 700 265
rect 635 235 645 255
rect 665 245 700 255
rect 665 235 675 245
rect 635 225 675 235
rect 485 210 550 220
rect 530 195 550 210
rect 230 145 240 185
rect 260 145 270 185
rect 230 135 270 145
rect 330 185 370 195
rect 330 145 340 185
rect 360 145 370 185
rect 330 135 370 145
rect 430 185 470 195
rect 430 145 440 185
rect 460 145 470 185
rect 430 135 470 145
rect 530 185 570 195
rect 530 145 540 185
rect 560 145 570 185
rect 530 135 570 145
rect 50 115 70 135
rect 430 115 450 135
rect 50 105 800 115
rect 50 95 770 105
rect 760 85 770 95
rect 790 85 800 105
rect 760 75 800 85
rect -160 55 70 75
rect -220 -40 -180 -30
rect -155 25 -115 35
rect -155 5 -145 25
rect -125 5 -115 25
rect -25 25 15 35
rect -25 15 -15 25
rect -155 -5 -115 5
rect -50 5 -15 15
rect 5 5 15 25
rect -50 -5 15 5
rect 50 20 70 55
rect 330 30 370 40
rect 50 0 250 20
rect -400 -330 -380 -40
rect -300 -85 -280 -40
rect -155 -85 -135 -5
rect -50 -20 -30 -5
rect 50 -20 70 0
rect 230 -20 250 0
rect 330 10 340 30
rect 360 10 370 30
rect -75 -30 -30 -20
rect -75 -70 -60 -30
rect -40 -70 -30 -30
rect -75 -80 -30 -70
rect 30 -30 70 -20
rect 30 -70 40 -30
rect 60 -70 70 -30
rect 30 -80 70 -70
rect 130 -30 170 -20
rect 130 -70 140 -30
rect 160 -70 170 -30
rect 130 -80 170 -70
rect 230 -30 270 -20
rect 230 -70 240 -30
rect 260 -70 270 -30
rect 230 -80 270 -70
rect 330 -30 370 10
rect 685 30 725 40
rect 685 10 695 30
rect 715 20 725 30
rect 715 10 750 20
rect 685 0 750 10
rect 730 -20 750 0
rect 330 -70 340 -30
rect 360 -70 370 -30
rect 330 -80 370 -70
rect 430 -30 470 -20
rect 430 -70 440 -30
rect 460 -70 470 -30
rect 430 -80 470 -70
rect 530 -30 570 -20
rect 530 -70 540 -30
rect 560 -70 570 -30
rect 530 -80 570 -70
rect 630 -30 670 -20
rect 630 -70 640 -30
rect 660 -70 670 -30
rect 630 -80 670 -70
rect 730 -30 770 -20
rect 730 -70 740 -30
rect 760 -70 770 -30
rect 730 -80 770 -70
rect -300 -105 -135 -85
rect 530 -100 550 -80
rect 530 -120 765 -100
rect -10 -140 30 -130
rect -10 -160 0 -140
rect 20 -160 30 -140
rect -265 -175 -225 -165
rect -265 -185 -255 -175
rect -290 -195 -255 -185
rect -235 -195 -225 -175
rect -165 -175 -125 -165
rect -165 -185 -155 -175
rect -290 -205 -225 -195
rect -190 -195 -155 -185
rect -135 -195 -125 -175
rect -190 -205 -125 -195
rect -10 -170 30 -160
rect -290 -225 -270 -205
rect -190 -225 -170 -205
rect -10 -225 10 -170
rect 145 -175 185 -165
rect 145 -195 155 -175
rect 175 -185 185 -175
rect 290 -175 330 -165
rect 175 -195 210 -185
rect 145 -205 210 -195
rect 190 -225 210 -205
rect 290 -195 300 -175
rect 320 -195 330 -175
rect -360 -235 -270 -225
rect -360 -275 -350 -235
rect -330 -275 -300 -235
rect -280 -275 -270 -235
rect -360 -285 -270 -275
rect -210 -235 -170 -225
rect -210 -275 -200 -235
rect -180 -275 -170 -235
rect -210 -285 -170 -275
rect -110 -235 -70 -225
rect -110 -275 -100 -235
rect -80 -275 -70 -235
rect -110 -285 -70 -275
rect -10 -235 30 -225
rect -10 -275 0 -235
rect 20 -275 30 -235
rect -10 -285 30 -275
rect 90 -235 130 -225
rect 90 -275 100 -235
rect 120 -275 130 -235
rect 90 -285 130 -275
rect 190 -235 230 -225
rect 190 -275 200 -235
rect 220 -275 230 -235
rect 190 -285 230 -275
rect 290 -235 330 -195
rect 645 -175 685 -165
rect 645 -195 655 -175
rect 675 -185 685 -175
rect 745 -175 765 -120
rect 745 -185 785 -175
rect 675 -195 710 -185
rect 645 -205 710 -195
rect 690 -225 710 -205
rect 745 -205 755 -185
rect 775 -205 785 -185
rect 745 -215 785 -205
rect 290 -275 300 -235
rect 320 -275 330 -235
rect 290 -285 330 -275
rect 390 -235 430 -225
rect 390 -275 400 -235
rect 420 -275 430 -235
rect 390 -285 430 -275
rect 490 -235 530 -225
rect 490 -275 500 -235
rect 520 -275 530 -235
rect 490 -285 530 -275
rect 590 -235 630 -225
rect 590 -275 600 -235
rect 620 -275 630 -235
rect 590 -285 630 -275
rect 690 -235 730 -225
rect 690 -275 700 -235
rect 720 -275 730 -235
rect 690 -285 730 -275
rect -190 -305 -170 -285
rect -10 -305 10 -285
rect -190 -325 -90 -305
rect -10 -325 210 -305
rect -625 -340 -285 -330
rect -625 -350 -315 -340
rect -325 -360 -315 -350
rect -295 -360 -285 -340
rect -325 -370 -285 -360
rect -265 -405 -225 -395
rect -265 -415 -255 -405
rect -290 -425 -255 -415
rect -235 -425 -225 -405
rect -290 -435 -225 -425
rect -290 -450 -270 -435
rect -110 -450 -90 -325
rect 90 -405 130 -395
rect 90 -425 100 -405
rect 120 -425 130 -405
rect -360 -460 -270 -450
rect -360 -500 -350 -460
rect -330 -500 -300 -460
rect -280 -500 -270 -460
rect -360 -510 -270 -500
rect -210 -460 -170 -450
rect -210 -500 -200 -460
rect -180 -500 -170 -460
rect -210 -510 -170 -500
rect -110 -460 -70 -450
rect -110 -500 -100 -460
rect -80 -500 -70 -460
rect -110 -510 -70 -500
rect -10 -460 30 -450
rect -10 -500 0 -460
rect 20 -500 30 -460
rect -10 -510 30 -500
rect 90 -460 130 -425
rect 90 -500 100 -460
rect 120 -500 130 -460
rect 90 -510 130 -500
rect 190 -450 210 -325
rect 490 -315 510 -285
rect 490 -335 800 -315
rect 490 -355 510 -335
rect 310 -375 470 -355
rect 310 -450 330 -375
rect 190 -460 230 -450
rect 190 -500 200 -460
rect 220 -500 230 -460
rect 190 -510 230 -500
rect 290 -460 330 -450
rect 290 -500 300 -460
rect 320 -500 330 -460
rect 290 -510 330 -500
rect 390 -405 430 -395
rect 390 -425 400 -405
rect 420 -425 430 -405
rect 390 -460 430 -425
rect 390 -500 400 -460
rect 420 -500 430 -460
rect 450 -450 470 -375
rect 490 -365 530 -355
rect 490 -385 500 -365
rect 520 -385 530 -365
rect 490 -395 530 -385
rect 550 -365 780 -355
rect 550 -375 750 -365
rect 550 -450 570 -375
rect 740 -385 750 -375
rect 770 -385 780 -365
rect 740 -395 780 -385
rect 645 -405 685 -395
rect 645 -425 655 -405
rect 675 -415 685 -405
rect 675 -425 710 -415
rect 645 -435 710 -425
rect 690 -450 710 -435
rect 450 -460 570 -450
rect 450 -470 500 -460
rect 390 -510 430 -500
rect 490 -500 500 -470
rect 520 -470 570 -460
rect 590 -460 630 -450
rect 520 -500 530 -470
rect 490 -510 530 -500
rect 590 -500 600 -460
rect 620 -500 630 -460
rect 590 -510 630 -500
rect 690 -460 730 -450
rect 690 -500 700 -460
rect 720 -500 730 -460
rect 690 -510 730 -500
rect 210 -525 230 -510
rect 590 -525 610 -510
rect 210 -530 275 -525
rect 545 -530 610 -525
rect 210 -535 610 -530
rect 210 -550 245 -535
rect 235 -555 245 -550
rect 265 -550 555 -535
rect 265 -555 275 -550
rect 235 -565 275 -555
rect 545 -555 555 -550
rect 575 -550 610 -535
rect 575 -555 585 -550
rect 545 -565 585 -555
<< viali >>
rect -610 -30 -590 500
rect -210 -30 -190 500
rect 40 495 60 535
rect 90 495 110 535
rect 290 495 310 535
rect 490 495 510 535
rect 690 495 710 535
rect 705 435 740 455
rect 40 320 60 360
rect 90 320 110 360
rect 290 320 310 360
rect 490 320 510 360
rect 690 320 710 360
rect 240 240 260 255
rect 240 220 260 240
rect -110 145 -90 185
rect -60 145 -40 185
rect 140 145 160 185
rect 340 145 360 185
rect 540 145 560 185
rect -60 -70 -40 -30
rect 140 -70 160 -30
rect 340 -70 360 -30
rect 440 -70 460 -30
rect 640 -70 660 -30
rect 740 -70 760 -30
rect -350 -275 -330 -235
rect -300 -275 -280 -235
rect -100 -275 -80 -235
rect 100 -275 120 -235
rect 300 -275 320 -235
rect 400 -275 420 -235
rect 600 -275 620 -235
rect 700 -275 720 -235
rect -350 -500 -330 -460
rect -300 -500 -280 -460
rect -200 -500 -180 -460
rect 0 -500 20 -460
rect 100 -500 120 -460
rect 700 -500 720 -460
<< metal1 >>
rect -625 585 -135 605
rect -150 545 -135 585
rect -150 535 725 545
rect -625 500 -180 510
rect -625 -30 -610 500
rect -590 -30 -210 500
rect -190 -30 -180 500
rect -625 -40 -180 -30
rect -150 495 40 535
rect 60 495 90 535
rect 110 495 290 535
rect 310 495 490 535
rect 510 495 690 535
rect 710 495 725 535
rect -150 485 725 495
rect -150 370 -135 485
rect 690 455 755 465
rect 690 435 705 455
rect 740 435 755 455
rect 690 425 755 435
rect -150 360 725 370
rect -150 320 40 360
rect 60 320 90 360
rect 110 320 290 360
rect 310 320 490 360
rect 510 320 690 360
rect 710 320 725 360
rect -150 310 725 320
rect -445 -450 -410 -40
rect -150 -225 -135 310
rect 740 280 755 425
rect 230 265 755 280
rect 230 255 270 265
rect 230 220 240 255
rect 260 220 270 255
rect 230 210 270 220
rect -120 185 570 195
rect -120 145 -110 185
rect -90 145 -60 185
rect -40 145 140 185
rect 160 145 340 185
rect 360 145 540 185
rect 560 145 570 185
rect -120 135 570 145
rect -70 -20 -30 135
rect 740 20 755 265
rect 740 0 800 20
rect -75 -30 775 -20
rect -75 -70 -60 -30
rect -40 -70 140 -30
rect 160 -70 340 -30
rect 360 -70 440 -30
rect 460 -70 640 -30
rect 660 -70 740 -30
rect 760 -70 775 -30
rect -75 -80 775 -70
rect -360 -235 735 -225
rect -360 -275 -350 -235
rect -330 -275 -300 -235
rect -280 -275 -100 -235
rect -80 -275 100 -235
rect 120 -275 300 -235
rect 320 -275 400 -235
rect 420 -275 600 -235
rect 620 -275 700 -235
rect 720 -275 735 -235
rect -360 -285 735 -275
rect 750 -450 765 -80
rect -445 -460 765 -450
rect -445 -500 -350 -460
rect -330 -500 -300 -460
rect -280 -500 -200 -460
rect -180 -500 0 -460
rect 20 -500 100 -460
rect 120 -500 700 -460
rect 720 -500 765 -460
rect -445 -510 765 -500
<< labels >>
rlabel metal1 -625 595 -625 595 7 VP
port 1 w
rlabel metal1 -625 235 -625 235 7 VN
port 2 w
rlabel locali -625 -340 -625 -340 7 Rbias
port 3 w
rlabel metal1 800 10 800 10 3 Vbn
port 4 e
rlabel locali 800 -325 800 -325 3 Vc
port 5 e
<< end >>
