* SPICE3 file created from dacladder.ext - technology: sky130A


* Top level circuit dacladder

X0 branch2 VP branch1 VN sky130_fd_pr__nfet_01v8 ad=1.425e+13p pd=6.2e+07u as=1.425e+13p ps=6.2e+07u w=5.7e+06u l=1.4e+06u
X1 VP VN VN VN sky130_fd_pr__nfet_01v8 ad=1.995e+13p pd=8.68e+07u as=1.653e+13p ps=7.42e+07u w=5.7e+06u l=1.4e+06u
X2 branch1 VP branch0 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.55e+12p ps=3.72e+07u w=5.7e+06u l=1.4e+06u
X3 branch3 VP branch2 VN sky130_fd_pr__nfet_01v8 ad=1.425e+13p pd=6.2e+07u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X4 branch4 VP branch3 VN sky130_fd_pr__nfet_01v8 ad=1.425e+13p pd=6.2e+07u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X5 branch6 VP branch5 VN sky130_fd_pr__nfet_01v8 ad=1.14e+13p pd=4.96e+07u as=1.425e+13p ps=6.2e+07u w=5.7e+06u l=1.4e+06u
X6 VN VN branch6 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X7 branch0 VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X8 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.7e+12p ps=2.48e+07u w=5.7e+06u l=1.4e+06u
X9 branch4 VP branch3 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X10 VP VP branch2 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X11 branch0 VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X12 VP VP branch4 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X13 branch5 VP branch4 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X14 Iout VP branch6 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X15 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X16 VP VP branch0 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X17 branch3 VP branch2 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X18 VP VP branch1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X19 branch5 VP branch4 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X20 VP VP branch3 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X21 Iout VP branch6 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X22 branch2 VP branch1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X23 branch6 VP branch5 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X24 VP VP branch5 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X25 branch1 VP branch0 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X26 branch0 VP VP VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
.end

