* SPICE3 file created from /home/jonah/VLSI/VLSI-MP4/design-files/layout/dac.ext - technology: sky130A

.subckt biasgen Vc Rbias Vbn VN VP
X0 a_50_260# a_50_n170# VP VP sky130_fd_pr__pfet_01v8 ad=3.5e+11p pd=2.4e+06u as=5.25e+12p ps=3.6e+07u w=700000u l=500000u
X1 VN VN a_50_260# VN sky130_fd_pr__nfet_01v8 ad=1.085e+13p pd=6.04e+07u as=7e+11p ps=4.8e+06u w=700000u l=500000u
X2 a_n30_n580# VN VN VN sky130_fd_pr__nfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X3 a_n430_n580# a_n430_n580# VP VP sky130_fd_pr__pfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X4 a_50_n170# VN VN VN sky130_fd_pr__nfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X5 VN a_n30_n580# a_570_n1030# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.05e+12p ps=7.2e+06u w=700000u l=500000u
X6 VP a_n430_n580# a_n430_n580# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X7 a_n1050_n90# VN VN VN sky130_fd_pr__nfet_01v8 ad=5.6e+12p pd=2.44e+07u as=0p ps=0u w=5.6e+06u l=500000u
X8 Rbias a_n1050_n90# a_n1050_n90# VN sky130_fd_pr__nfet_01v8 ad=2.8e+12p pd=1.22e+07u as=0p ps=0u w=5.6e+06u l=500000u
X9 a_50_n170# VP VP VP sky130_fd_pr__pfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X10 a_50_260# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X11 a_570_n1030# a_n30_n580# a_n30_n580# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X12 a_n1050_n90# a_50_260# VP VP sky130_fd_pr__pfet_01v8 ad=7e+11p pd=4.8e+06u as=0p ps=0u w=700000u l=500000u
X13 VN Vbn Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5e+11p ps=2.4e+06u w=700000u l=500000u
X14 VN VN a_50_n170# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X15 VP a_50_260# Vbn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.5e+11p ps=2.4e+06u w=700000u l=500000u
X16 Vc Vc a_570_n1030# VN sky130_fd_pr__nfet_01v8 ad=3.5e+11p pd=2.4e+06u as=0p ps=0u w=700000u l=500000u
X17 Vc a_50_260# VP VP sky130_fd_pr__pfet_01v8 ad=3.5e+11p pd=2.4e+06u as=0p ps=0u w=700000u l=500000u
X18 VN Rbias a_n430_n580# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5e+11p ps=2.4e+06u w=700000u l=500000u
X19 VN VN a_n1050_n90# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.6e+06u l=500000u
X20 a_570_n1030# Vc Vc VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X21 VN Vbn a_50_260# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X22 a_n30_n580# a_n430_n580# VP VP sky130_fd_pr__pfet_01v8 ad=3.5e+11p pd=2.4e+06u as=0p ps=0u w=700000u l=500000u
X23 a_n430_n580# Rbias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X24 VP a_50_260# a_n1050_n90# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X25 a_50_n170# a_50_n170# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X26 VP a_50_n170# a_50_260# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X27 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X28 a_50_n170# a_n1050_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X29 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X30 VP a_n430_n580# a_n30_n580# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X31 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X32 VP a_50_n170# a_50_n170# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X33 VP VP a_n1050_n90# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X34 a_50_260# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X35 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X36 a_570_n1030# a_n30_n580# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X37 VP a_50_260# Vc VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X38 VN a_n1050_n90# a_50_n170# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X39 a_n1050_n90# a_n1050_n90# Rbias VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.6e+06u l=500000u
X40 Vbn Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X41 a_n30_n580# a_n30_n580# a_570_n1030# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X42 Vbn a_50_260# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X43 VP VP a_50_n170# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X44 VP VP a_n430_n580# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X45 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X46 a_n430_n580# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X47 VN VN a_n30_n580# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X48 a_n1050_n90# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X49 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
.ends

.subckt dacladder Iout branch0 branch1 branch2 branch3 branch4 branch5 branch6 VN
+ VP
X0 branch2 VP branch1 VN sky130_fd_pr__nfet_01v8 ad=1.425e+13p pd=6.2e+07u as=1.425e+13p ps=6.2e+07u w=5.7e+06u l=1.4e+06u
X1 VP VN VN VN sky130_fd_pr__nfet_01v8 ad=1.995e+13p pd=8.68e+07u as=1.653e+13p ps=7.42e+07u w=5.7e+06u l=1.4e+06u
X2 branch1 VP branch0 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.55e+12p ps=3.72e+07u w=5.7e+06u l=1.4e+06u
X3 branch3 VP branch2 VN sky130_fd_pr__nfet_01v8 ad=1.425e+13p pd=6.2e+07u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X4 branch4 VP branch3 VN sky130_fd_pr__nfet_01v8 ad=1.425e+13p pd=6.2e+07u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X5 branch6 VP branch5 VN sky130_fd_pr__nfet_01v8 ad=1.14e+13p pd=4.96e+07u as=1.425e+13p ps=6.2e+07u w=5.7e+06u l=1.4e+06u
X6 VN VN branch6 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X7 branch0 VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X8 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.7e+12p ps=2.48e+07u w=5.7e+06u l=1.4e+06u
X9 branch4 VP branch3 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X10 VP VP branch2 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X11 branch0 VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X12 VP VP branch4 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X13 branch5 VP branch4 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X14 Iout VP branch6 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X15 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X16 VP VP branch0 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X17 branch3 VP branch2 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X18 VP VP branch1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X19 branch5 VP branch4 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X20 VP VP branch3 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X21 Iout VP branch6 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X22 branch2 VP branch1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X23 branch6 VP branch5 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X24 VP VP branch5 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X25 branch1 VP branch0 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
X26 branch0 VP VP VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.7e+06u l=1.4e+06u
.ends

.subckt branchl Vc branch0 branch1 Vbn branch2 branch3 branch4 branch5 branch6 VN
+ VP
X0 a_2390_n90# a_2370_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=1.5925e+13p ps=7.77e+07u w=3.15e+06u l=300000u
X1 a_4700_720# a_3710_n90# VN VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=0p ps=0u w=1.4e+06u l=500000u
X2 a_n250_n90# a_n270_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X3 VN b5in a_6330_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X4 VP b6in a_7650_650# VP sky130_fd_pr__pfet_01v8 ad=1.1025e+13p pd=5.11e+07u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X5 a_2060_720# a_1070_n90# VN VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=0p ps=0u w=1.4e+06u l=500000u
X6 a_7670_n90# a_7650_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=1.1025e+13p ps=5.11e+07u w=3.15e+06u l=300000u
X7 VN b3in a_3690_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X8 a_3710_n90# b3in Vbn VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=1.1025e+13p ps=5.11e+07u w=3.15e+06u l=300000u
X9 a_8660_720# Vc branch6 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X10 a_6350_n90# a_6330_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X11 VP b5in a_6330_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X12 a_n250_n90# b0in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X13 VN b2in a_2370_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X14 a_740_720# Vc branch0 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X15 a_3710_n90# a_3690_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X16 a_2390_n90# b2in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X17 a_6350_n90# a_6330_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X18 a_8660_720# a_7670_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X19 a_7340_720# Vc branch5 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X20 a_5030_n90# a_5010_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X21 VP b4in a_5010_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X22 VP b2in a_2370_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X23 a_740_720# a_n250_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X24 VN b1in a_1050_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X25 a_2390_n90# a_2370_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X26 a_1070_n90# b1in Vbn VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X27 a_5030_n90# a_5010_650# VN VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X28 a_7340_720# a_6350_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X29 a_n250_n90# a_n270_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X30 VP b3in a_3690_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X31 a_3380_720# Vc branch2 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X32 VP b1in a_1050_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X33 a_1070_n90# a_1050_650# Vbn VP sky130_fd_pr__pfet_01v8 ad=1.575e+12p pd=7.3e+06u as=0p ps=0u w=3.15e+06u l=300000u
X34 a_3710_n90# a_3690_650# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X35 a_6350_n90# b5in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X36 a_1070_n90# a_1050_650# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X37 a_3380_720# a_2390_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X38 VN b0in a_n270_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X39 a_6020_720# Vc branch4 VN sky130_fd_pr__nfet_01v8 ad=1.4e+12p pd=7.6e+06u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X40 VN b4in a_5010_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X41 VP b0in a_n270_650# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X42 a_6020_720# a_5030_n90# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=500000u
X43 a_4700_720# Vc branch3 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X44 a_7670_n90# b6in Vbn VN sky130_fd_pr__nfet_01v8 ad=3.15e+12p pd=1.46e+07u as=0p ps=0u w=3.15e+06u l=300000u
X45 VN b6in a_7650_650# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.575e+12p ps=7.3e+06u w=3.15e+06u l=300000u
X46 a_7670_n90# a_7650_650# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
X47 a_2060_720# Vc branch1 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7e+11p ps=3.8e+06u w=1.4e+06u l=500000u
X48 a_5030_n90# b4in Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.15e+06u l=300000u
.ends


* Top level circuit /home/jonah/VLSI/VLSI-MP4/design-files/layout/dac

Xbiasgen_0 branchl_0/Vc Rbias branchl_0/Vbn VN VP biasgen
Xdacladder_0 Iout branchl_0/branch0 branchl_0/branch1 branchl_0/branch2 branchl_0/branch3
+ branchl_0/branch4 branchl_0/branch5 branchl_0/branch6 VN VP dacladder
Xbranchl_0 branchl_0/Vc branchl_0/branch0 branchl_0/branch1 branchl_0/Vbn branchl_0/branch2
+ branchl_0/branch3 branchl_0/branch4 branchl_0/branch5 branchl_0/branch6 VN VP branchl
.end

