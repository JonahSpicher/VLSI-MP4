magic
tech sky130A
timestamp 1617823527
<< nwell >>
rect -205 320 175 675
rect 455 320 835 675
rect 1115 320 1495 675
rect 1775 320 2155 675
rect 2435 320 2815 675
rect 3095 320 3475 675
rect 3755 320 4135 675
<< nmos >>
rect 320 360 370 500
rect 980 360 1030 500
rect 1640 360 1690 500
rect 2300 360 2350 500
rect 2960 360 3010 500
rect 3620 360 3670 500
rect 4280 360 4330 500
rect -155 -45 -125 270
rect 5 -45 35 270
rect 85 -45 115 270
rect 325 130 375 270
rect 505 -45 535 270
rect 665 -45 695 270
rect 745 -45 775 270
rect 985 130 1035 270
rect 1165 -45 1195 270
rect 1325 -45 1355 270
rect 1405 -45 1435 270
rect 1645 130 1695 270
rect 1825 -45 1855 270
rect 1985 -45 2015 270
rect 2065 -45 2095 270
rect 2305 130 2355 270
rect 2485 -45 2515 270
rect 2645 -45 2675 270
rect 2725 -45 2755 270
rect 2965 130 3015 270
rect 3145 -45 3175 270
rect 3305 -45 3335 270
rect 3385 -45 3415 270
rect 3625 130 3675 270
rect 3805 -45 3835 270
rect 3965 -45 3995 270
rect 4045 -45 4075 270
rect 4285 130 4335 270
<< pmos >>
rect -135 340 -105 655
rect 25 340 55 655
rect 525 340 555 655
rect 685 340 715 655
rect 1185 340 1215 655
rect 1345 340 1375 655
rect 1845 340 1875 655
rect 2005 340 2035 655
rect 2505 340 2535 655
rect 2665 340 2695 655
rect 3165 340 3195 655
rect 3325 340 3355 655
rect 3825 340 3855 655
rect 3985 340 4015 655
<< ndiff >>
rect 270 485 320 500
rect 270 375 285 485
rect 305 375 320 485
rect 270 360 320 375
rect 370 485 420 500
rect 370 375 385 485
rect 405 375 420 485
rect 370 360 420 375
rect 930 485 980 500
rect 930 375 945 485
rect 965 375 980 485
rect 930 360 980 375
rect 1030 485 1080 500
rect 1030 375 1045 485
rect 1065 375 1080 485
rect 1030 360 1080 375
rect 1590 485 1640 500
rect 1590 375 1605 485
rect 1625 375 1640 485
rect 1590 360 1640 375
rect 1690 485 1740 500
rect 1690 375 1705 485
rect 1725 375 1740 485
rect 1690 360 1740 375
rect 2250 485 2300 500
rect 2250 375 2265 485
rect 2285 375 2300 485
rect 2250 360 2300 375
rect 2350 485 2400 500
rect 2350 375 2365 485
rect 2385 375 2400 485
rect 2350 360 2400 375
rect 2910 485 2960 500
rect 2910 375 2925 485
rect 2945 375 2960 485
rect 2910 360 2960 375
rect 3010 485 3060 500
rect 3010 375 3025 485
rect 3045 375 3060 485
rect 3010 360 3060 375
rect 3570 485 3620 500
rect 3570 375 3585 485
rect 3605 375 3620 485
rect 3570 360 3620 375
rect 3670 485 3720 500
rect 3670 375 3685 485
rect 3705 375 3720 485
rect 3670 360 3720 375
rect 4230 485 4280 500
rect 4230 375 4245 485
rect 4265 375 4280 485
rect 4230 360 4280 375
rect 4330 485 4380 500
rect 4330 375 4345 485
rect 4365 375 4380 485
rect 4330 360 4380 375
rect -205 255 -155 270
rect -205 -30 -190 255
rect -170 -30 -155 255
rect -205 -45 -155 -30
rect -125 255 -75 270
rect -125 -30 -110 255
rect -90 -30 -75 255
rect -125 -45 -75 -30
rect -45 255 5 270
rect -45 -30 -30 255
rect -10 -30 5 255
rect -45 -45 5 -30
rect 35 255 85 270
rect 35 -30 50 255
rect 70 -30 85 255
rect 35 -45 85 -30
rect 115 255 165 270
rect 115 -30 130 255
rect 150 -30 165 255
rect 115 -45 165 -30
rect 275 255 325 270
rect 275 145 290 255
rect 310 145 325 255
rect 275 130 325 145
rect 375 255 425 270
rect 375 145 390 255
rect 410 145 425 255
rect 375 130 425 145
rect 455 255 505 270
rect 455 -30 470 255
rect 490 -30 505 255
rect 455 -45 505 -30
rect 535 255 585 270
rect 535 -30 550 255
rect 570 -30 585 255
rect 535 -45 585 -30
rect 615 255 665 270
rect 615 -30 630 255
rect 650 -30 665 255
rect 615 -45 665 -30
rect 695 255 745 270
rect 695 -30 710 255
rect 730 -30 745 255
rect 695 -45 745 -30
rect 775 255 825 270
rect 775 -30 790 255
rect 810 -30 825 255
rect 775 -45 825 -30
rect 935 255 985 270
rect 935 145 950 255
rect 970 145 985 255
rect 935 130 985 145
rect 1035 255 1085 270
rect 1035 145 1050 255
rect 1070 145 1085 255
rect 1035 130 1085 145
rect 1115 255 1165 270
rect 1115 -30 1130 255
rect 1150 -30 1165 255
rect 1115 -45 1165 -30
rect 1195 255 1245 270
rect 1195 -30 1210 255
rect 1230 -30 1245 255
rect 1195 -45 1245 -30
rect 1275 255 1325 270
rect 1275 -30 1290 255
rect 1310 -30 1325 255
rect 1275 -45 1325 -30
rect 1355 255 1405 270
rect 1355 -30 1370 255
rect 1390 -30 1405 255
rect 1355 -45 1405 -30
rect 1435 255 1485 270
rect 1435 -30 1450 255
rect 1470 -30 1485 255
rect 1435 -45 1485 -30
rect 1595 255 1645 270
rect 1595 145 1610 255
rect 1630 145 1645 255
rect 1595 130 1645 145
rect 1695 255 1745 270
rect 1695 145 1710 255
rect 1730 145 1745 255
rect 1695 130 1745 145
rect 1775 255 1825 270
rect 1775 -30 1790 255
rect 1810 -30 1825 255
rect 1775 -45 1825 -30
rect 1855 255 1905 270
rect 1855 -30 1870 255
rect 1890 -30 1905 255
rect 1855 -45 1905 -30
rect 1935 255 1985 270
rect 1935 -30 1950 255
rect 1970 -30 1985 255
rect 1935 -45 1985 -30
rect 2015 255 2065 270
rect 2015 -30 2030 255
rect 2050 -30 2065 255
rect 2015 -45 2065 -30
rect 2095 255 2145 270
rect 2095 -30 2110 255
rect 2130 -30 2145 255
rect 2095 -45 2145 -30
rect 2255 255 2305 270
rect 2255 145 2270 255
rect 2290 145 2305 255
rect 2255 130 2305 145
rect 2355 255 2405 270
rect 2355 145 2370 255
rect 2390 145 2405 255
rect 2355 130 2405 145
rect 2435 255 2485 270
rect 2435 -30 2450 255
rect 2470 -30 2485 255
rect 2435 -45 2485 -30
rect 2515 255 2565 270
rect 2515 -30 2530 255
rect 2550 -30 2565 255
rect 2515 -45 2565 -30
rect 2595 255 2645 270
rect 2595 -30 2610 255
rect 2630 -30 2645 255
rect 2595 -45 2645 -30
rect 2675 255 2725 270
rect 2675 -30 2690 255
rect 2710 -30 2725 255
rect 2675 -45 2725 -30
rect 2755 255 2805 270
rect 2755 -30 2770 255
rect 2790 -30 2805 255
rect 2755 -45 2805 -30
rect 2915 255 2965 270
rect 2915 145 2930 255
rect 2950 145 2965 255
rect 2915 130 2965 145
rect 3015 255 3065 270
rect 3015 145 3030 255
rect 3050 145 3065 255
rect 3015 130 3065 145
rect 3095 255 3145 270
rect 3095 -30 3110 255
rect 3130 -30 3145 255
rect 3095 -45 3145 -30
rect 3175 255 3225 270
rect 3175 -30 3190 255
rect 3210 -30 3225 255
rect 3175 -45 3225 -30
rect 3255 255 3305 270
rect 3255 -30 3270 255
rect 3290 -30 3305 255
rect 3255 -45 3305 -30
rect 3335 255 3385 270
rect 3335 -30 3350 255
rect 3370 -30 3385 255
rect 3335 -45 3385 -30
rect 3415 255 3465 270
rect 3415 -30 3430 255
rect 3450 -30 3465 255
rect 3415 -45 3465 -30
rect 3575 255 3625 270
rect 3575 145 3590 255
rect 3610 145 3625 255
rect 3575 130 3625 145
rect 3675 255 3725 270
rect 3675 145 3690 255
rect 3710 145 3725 255
rect 3675 130 3725 145
rect 3755 255 3805 270
rect 3755 -30 3770 255
rect 3790 -30 3805 255
rect 3755 -45 3805 -30
rect 3835 255 3885 270
rect 3835 -30 3850 255
rect 3870 -30 3885 255
rect 3835 -45 3885 -30
rect 3915 255 3965 270
rect 3915 -30 3930 255
rect 3950 -30 3965 255
rect 3915 -45 3965 -30
rect 3995 255 4045 270
rect 3995 -30 4010 255
rect 4030 -30 4045 255
rect 3995 -45 4045 -30
rect 4075 255 4125 270
rect 4075 -30 4090 255
rect 4110 -30 4125 255
rect 4075 -45 4125 -30
rect 4235 255 4285 270
rect 4235 145 4250 255
rect 4270 145 4285 255
rect 4235 130 4285 145
rect 4335 255 4385 270
rect 4335 145 4350 255
rect 4370 145 4385 255
rect 4335 130 4385 145
<< pdiff >>
rect -185 640 -135 655
rect -185 355 -170 640
rect -150 355 -135 640
rect -185 340 -135 355
rect -105 640 -55 655
rect -105 355 -90 640
rect -70 355 -55 640
rect -105 340 -55 355
rect -25 640 25 655
rect -25 355 -10 640
rect 10 355 25 640
rect -25 340 25 355
rect 55 640 105 655
rect 55 355 70 640
rect 90 355 105 640
rect 475 640 525 655
rect 55 340 105 355
rect 475 355 490 640
rect 510 355 525 640
rect 475 340 525 355
rect 555 640 605 655
rect 555 355 570 640
rect 590 355 605 640
rect 555 340 605 355
rect 635 640 685 655
rect 635 355 650 640
rect 670 355 685 640
rect 635 340 685 355
rect 715 640 765 655
rect 715 355 730 640
rect 750 355 765 640
rect 1135 640 1185 655
rect 715 340 765 355
rect 1135 355 1150 640
rect 1170 355 1185 640
rect 1135 340 1185 355
rect 1215 640 1265 655
rect 1215 355 1230 640
rect 1250 355 1265 640
rect 1215 340 1265 355
rect 1295 640 1345 655
rect 1295 355 1310 640
rect 1330 355 1345 640
rect 1295 340 1345 355
rect 1375 640 1425 655
rect 1375 355 1390 640
rect 1410 355 1425 640
rect 1795 640 1845 655
rect 1375 340 1425 355
rect 1795 355 1810 640
rect 1830 355 1845 640
rect 1795 340 1845 355
rect 1875 640 1925 655
rect 1875 355 1890 640
rect 1910 355 1925 640
rect 1875 340 1925 355
rect 1955 640 2005 655
rect 1955 355 1970 640
rect 1990 355 2005 640
rect 1955 340 2005 355
rect 2035 640 2085 655
rect 2035 355 2050 640
rect 2070 355 2085 640
rect 2455 640 2505 655
rect 2035 340 2085 355
rect 2455 355 2470 640
rect 2490 355 2505 640
rect 2455 340 2505 355
rect 2535 640 2585 655
rect 2535 355 2550 640
rect 2570 355 2585 640
rect 2535 340 2585 355
rect 2615 640 2665 655
rect 2615 355 2630 640
rect 2650 355 2665 640
rect 2615 340 2665 355
rect 2695 640 2745 655
rect 2695 355 2710 640
rect 2730 355 2745 640
rect 3115 640 3165 655
rect 2695 340 2745 355
rect 3115 355 3130 640
rect 3150 355 3165 640
rect 3115 340 3165 355
rect 3195 640 3245 655
rect 3195 355 3210 640
rect 3230 355 3245 640
rect 3195 340 3245 355
rect 3275 640 3325 655
rect 3275 355 3290 640
rect 3310 355 3325 640
rect 3275 340 3325 355
rect 3355 640 3405 655
rect 3355 355 3370 640
rect 3390 355 3405 640
rect 3775 640 3825 655
rect 3355 340 3405 355
rect 3775 355 3790 640
rect 3810 355 3825 640
rect 3775 340 3825 355
rect 3855 640 3905 655
rect 3855 355 3870 640
rect 3890 355 3905 640
rect 3855 340 3905 355
rect 3935 640 3985 655
rect 3935 355 3950 640
rect 3970 355 3985 640
rect 3935 340 3985 355
rect 4015 640 4065 655
rect 4015 355 4030 640
rect 4050 355 4065 640
rect 4015 340 4065 355
<< ndiffc >>
rect 285 375 305 485
rect 385 375 405 485
rect 945 375 965 485
rect 1045 375 1065 485
rect 1605 375 1625 485
rect 1705 375 1725 485
rect 2265 375 2285 485
rect 2365 375 2385 485
rect 2925 375 2945 485
rect 3025 375 3045 485
rect 3585 375 3605 485
rect 3685 375 3705 485
rect 4245 375 4265 485
rect 4345 375 4365 485
rect -190 -30 -170 255
rect -110 -30 -90 255
rect -30 -30 -10 255
rect 50 -30 70 255
rect 130 -30 150 255
rect 290 145 310 255
rect 390 145 410 255
rect 470 -30 490 255
rect 550 -30 570 255
rect 630 -30 650 255
rect 710 -30 730 255
rect 790 -30 810 255
rect 950 145 970 255
rect 1050 145 1070 255
rect 1130 -30 1150 255
rect 1210 -30 1230 255
rect 1290 -30 1310 255
rect 1370 -30 1390 255
rect 1450 -30 1470 255
rect 1610 145 1630 255
rect 1710 145 1730 255
rect 1790 -30 1810 255
rect 1870 -30 1890 255
rect 1950 -30 1970 255
rect 2030 -30 2050 255
rect 2110 -30 2130 255
rect 2270 145 2290 255
rect 2370 145 2390 255
rect 2450 -30 2470 255
rect 2530 -30 2550 255
rect 2610 -30 2630 255
rect 2690 -30 2710 255
rect 2770 -30 2790 255
rect 2930 145 2950 255
rect 3030 145 3050 255
rect 3110 -30 3130 255
rect 3190 -30 3210 255
rect 3270 -30 3290 255
rect 3350 -30 3370 255
rect 3430 -30 3450 255
rect 3590 145 3610 255
rect 3690 145 3710 255
rect 3770 -30 3790 255
rect 3850 -30 3870 255
rect 3930 -30 3950 255
rect 4010 -30 4030 255
rect 4090 -30 4110 255
rect 4250 145 4270 255
rect 4350 145 4370 255
<< pdiffc >>
rect -170 355 -150 640
rect -90 355 -70 640
rect -10 355 10 640
rect 70 355 90 640
rect 490 355 510 640
rect 570 355 590 640
rect 650 355 670 640
rect 730 355 750 640
rect 1150 355 1170 640
rect 1230 355 1250 640
rect 1310 355 1330 640
rect 1390 355 1410 640
rect 1810 355 1830 640
rect 1890 355 1910 640
rect 1970 355 1990 640
rect 2050 355 2070 640
rect 2470 355 2490 640
rect 2550 355 2570 640
rect 2630 355 2650 640
rect 2710 355 2730 640
rect 3130 355 3150 640
rect 3210 355 3230 640
rect 3290 355 3310 640
rect 3370 355 3390 640
rect 3790 355 3810 640
rect 3870 355 3890 640
rect 3950 355 3970 640
rect 4030 355 4050 640
<< psubdiff >>
rect 195 255 245 270
rect 195 -30 210 255
rect 230 -30 245 255
rect 195 -45 245 -30
rect 855 255 905 270
rect 855 -30 870 255
rect 890 -30 905 255
rect 855 -45 905 -30
rect 1515 255 1565 270
rect 1515 -30 1530 255
rect 1550 -30 1565 255
rect 1515 -45 1565 -30
rect 2175 255 2225 270
rect 2175 -30 2190 255
rect 2210 -30 2225 255
rect 2175 -45 2225 -30
rect 2835 255 2885 270
rect 2835 -30 2850 255
rect 2870 -30 2885 255
rect 2835 -45 2885 -30
rect 3495 255 3545 270
rect 3495 -30 3510 255
rect 3530 -30 3545 255
rect 3495 -45 3545 -30
rect 4155 255 4205 270
rect 4155 -30 4170 255
rect 4190 -30 4205 255
rect 4155 -45 4205 -30
<< nsubdiff >>
rect 105 640 155 655
rect 105 355 120 640
rect 140 355 155 640
rect 105 340 155 355
rect 765 640 815 655
rect 765 355 780 640
rect 800 355 815 640
rect 765 340 815 355
rect 1425 640 1475 655
rect 1425 355 1440 640
rect 1460 355 1475 640
rect 1425 340 1475 355
rect 2085 640 2135 655
rect 2085 355 2100 640
rect 2120 355 2135 640
rect 2085 340 2135 355
rect 2745 640 2795 655
rect 2745 355 2760 640
rect 2780 355 2795 640
rect 2745 340 2795 355
rect 3405 640 3455 655
rect 3405 355 3420 640
rect 3440 355 3455 640
rect 3405 340 3455 355
rect 4065 640 4115 655
rect 4065 355 4080 640
rect 4100 355 4115 640
rect 4065 340 4115 355
<< psubdiffcont >>
rect 210 -30 230 255
rect 870 -30 890 255
rect 1530 -30 1550 255
rect 2190 -30 2210 255
rect 2850 -30 2870 255
rect 3510 -30 3530 255
rect 4170 -30 4190 255
<< nsubdiffcont >>
rect 120 355 140 640
rect 780 355 800 640
rect 1440 355 1460 640
rect 2100 355 2120 640
rect 2760 355 2780 640
rect 3420 355 3440 640
rect 4080 355 4100 640
<< poly >>
rect -135 700 -95 710
rect -135 680 -125 700
rect -105 680 -95 700
rect -135 670 -95 680
rect 525 700 565 710
rect 525 680 535 700
rect 555 680 565 700
rect 525 670 565 680
rect 1185 700 1225 710
rect 1185 680 1195 700
rect 1215 680 1225 700
rect 1185 670 1225 680
rect 1845 700 1885 710
rect 1845 680 1855 700
rect 1875 680 1885 700
rect 1845 670 1885 680
rect 2505 700 2545 710
rect 2505 680 2515 700
rect 2535 680 2545 700
rect 2505 670 2545 680
rect 3165 700 3205 710
rect 3165 680 3175 700
rect 3195 680 3205 700
rect 3165 670 3205 680
rect 3825 700 3865 710
rect 3825 680 3835 700
rect 3855 680 3865 700
rect 3825 670 3865 680
rect -135 655 -105 670
rect 25 655 55 670
rect 525 655 555 670
rect 685 655 715 670
rect 1185 655 1215 670
rect 1345 655 1375 670
rect 1845 655 1875 670
rect 2005 655 2035 670
rect 2505 655 2535 670
rect 2665 655 2695 670
rect 3165 655 3195 670
rect 3325 655 3355 670
rect 3825 655 3855 670
rect 3985 655 4015 670
rect 330 545 370 555
rect 330 525 340 545
rect 360 525 370 545
rect 330 515 370 525
rect 320 500 370 515
rect 320 345 370 360
rect 990 545 1030 555
rect 990 525 1000 545
rect 1020 525 1030 545
rect 990 515 1030 525
rect 980 500 1030 515
rect 980 345 1030 360
rect 1650 545 1690 555
rect 1650 525 1660 545
rect 1680 525 1690 545
rect 1650 515 1690 525
rect 1640 500 1690 515
rect 1640 345 1690 360
rect 2310 545 2350 555
rect 2310 525 2320 545
rect 2340 525 2350 545
rect 2310 515 2350 525
rect 2300 500 2350 515
rect 2300 345 2350 360
rect 2970 545 3010 555
rect 2970 525 2980 545
rect 3000 525 3010 545
rect 2970 515 3010 525
rect 2960 500 3010 515
rect 2960 345 3010 360
rect 3630 545 3670 555
rect 3630 525 3640 545
rect 3660 525 3670 545
rect 3630 515 3670 525
rect 3620 500 3670 515
rect 3620 345 3670 360
rect 4290 545 4330 555
rect 4290 525 4300 545
rect 4320 525 4330 545
rect 4290 515 4330 525
rect 4280 500 4330 515
rect 4280 345 4330 360
rect -135 325 -105 340
rect 25 330 55 340
rect 5 315 55 330
rect 525 325 555 340
rect 685 330 715 340
rect 80 315 120 325
rect -155 270 -125 285
rect 5 270 35 315
rect 80 295 90 315
rect 110 295 120 315
rect 80 285 120 295
rect 260 315 300 325
rect 260 295 270 315
rect 290 300 300 315
rect 665 315 715 330
rect 1185 325 1215 340
rect 1345 330 1375 340
rect 740 315 780 325
rect 290 295 340 300
rect 260 285 340 295
rect 85 270 115 285
rect 325 270 375 285
rect 505 270 535 285
rect 665 270 695 315
rect 740 295 750 315
rect 770 295 780 315
rect 740 285 780 295
rect 920 315 960 325
rect 920 295 930 315
rect 950 300 960 315
rect 1325 315 1375 330
rect 1845 325 1875 340
rect 2005 330 2035 340
rect 1400 315 1440 325
rect 950 295 1000 300
rect 920 285 1000 295
rect 745 270 775 285
rect 985 270 1035 285
rect 1165 270 1195 285
rect 1325 270 1355 315
rect 1400 295 1410 315
rect 1430 295 1440 315
rect 1400 285 1440 295
rect 1580 315 1620 325
rect 1580 295 1590 315
rect 1610 300 1620 315
rect 1985 315 2035 330
rect 2505 325 2535 340
rect 2665 330 2695 340
rect 2060 315 2100 325
rect 1610 295 1660 300
rect 1580 285 1660 295
rect 1405 270 1435 285
rect 1645 270 1695 285
rect 1825 270 1855 285
rect 1985 270 2015 315
rect 2060 295 2070 315
rect 2090 295 2100 315
rect 2060 285 2100 295
rect 2240 315 2280 325
rect 2240 295 2250 315
rect 2270 300 2280 315
rect 2645 315 2695 330
rect 3165 325 3195 340
rect 3325 330 3355 340
rect 2720 315 2760 325
rect 2270 295 2320 300
rect 2240 285 2320 295
rect 2065 270 2095 285
rect 2305 270 2355 285
rect 2485 270 2515 285
rect 2645 270 2675 315
rect 2720 295 2730 315
rect 2750 295 2760 315
rect 2720 285 2760 295
rect 2900 315 2940 325
rect 2900 295 2910 315
rect 2930 300 2940 315
rect 3305 315 3355 330
rect 3825 325 3855 340
rect 3985 330 4015 340
rect 3380 315 3420 325
rect 2930 295 2980 300
rect 2900 285 2980 295
rect 2725 270 2755 285
rect 2965 270 3015 285
rect 3145 270 3175 285
rect 3305 270 3335 315
rect 3380 295 3390 315
rect 3410 295 3420 315
rect 3380 285 3420 295
rect 3560 315 3600 325
rect 3560 295 3570 315
rect 3590 300 3600 315
rect 3965 315 4015 330
rect 4040 315 4080 325
rect 3590 295 3640 300
rect 3560 285 3640 295
rect 3385 270 3415 285
rect 3625 270 3675 285
rect 3805 270 3835 285
rect 3965 270 3995 315
rect 4040 295 4050 315
rect 4070 295 4080 315
rect 4040 285 4080 295
rect 4220 315 4260 325
rect 4220 295 4230 315
rect 4250 300 4260 315
rect 4250 295 4300 300
rect 4220 285 4300 295
rect 4045 270 4075 285
rect 4285 270 4335 285
rect 325 115 375 130
rect 985 115 1035 130
rect 1645 115 1695 130
rect 2305 115 2355 130
rect 2965 115 3015 130
rect 3625 115 3675 130
rect 4285 115 4335 130
rect -155 -55 -125 -45
rect 5 -55 35 -45
rect -155 -70 35 -55
rect 85 -60 115 -45
rect 505 -55 535 -45
rect 665 -55 695 -45
rect 505 -70 695 -55
rect 745 -60 775 -45
rect 1165 -55 1195 -45
rect 1325 -55 1355 -45
rect 1165 -70 1355 -55
rect 1405 -60 1435 -45
rect 1825 -55 1855 -45
rect 1985 -55 2015 -45
rect 1825 -70 2015 -55
rect 2065 -60 2095 -45
rect 2485 -55 2515 -45
rect 2645 -55 2675 -45
rect 2485 -70 2675 -55
rect 2725 -60 2755 -45
rect 3145 -55 3175 -45
rect 3305 -55 3335 -45
rect 3145 -70 3335 -55
rect 3385 -60 3415 -45
rect 3805 -55 3835 -45
rect 3965 -55 3995 -45
rect 3805 -70 3995 -55
rect 4045 -60 4075 -45
rect -155 -75 -115 -70
rect -155 -95 -145 -75
rect -125 -95 -115 -75
rect -155 -105 -115 -95
rect 505 -75 545 -70
rect 505 -95 515 -75
rect 535 -95 545 -75
rect 505 -105 545 -95
rect 1165 -75 1205 -70
rect 1165 -95 1175 -75
rect 1195 -95 1205 -75
rect 1165 -105 1205 -95
rect 1825 -75 1865 -70
rect 1825 -95 1835 -75
rect 1855 -95 1865 -75
rect 1825 -105 1865 -95
rect 2485 -75 2525 -70
rect 2485 -95 2495 -75
rect 2515 -95 2525 -75
rect 2485 -105 2525 -95
rect 3145 -75 3185 -70
rect 3145 -95 3155 -75
rect 3175 -95 3185 -75
rect 3145 -105 3185 -95
rect 3805 -75 3845 -70
rect 3805 -95 3815 -75
rect 3835 -95 3845 -75
rect 3805 -105 3845 -95
<< polycont >>
rect -125 680 -105 700
rect 535 680 555 700
rect 1195 680 1215 700
rect 1855 680 1875 700
rect 2515 680 2535 700
rect 3175 680 3195 700
rect 3835 680 3855 700
rect 340 525 360 545
rect 1000 525 1020 545
rect 1660 525 1680 545
rect 2320 525 2340 545
rect 2980 525 3000 545
rect 3640 525 3660 545
rect 4300 525 4320 545
rect 90 295 110 315
rect 270 295 290 315
rect 750 295 770 315
rect 930 295 950 315
rect 1410 295 1430 315
rect 1590 295 1610 315
rect 2070 295 2090 315
rect 2250 295 2270 315
rect 2730 295 2750 315
rect 2910 295 2930 315
rect 3390 295 3410 315
rect 3570 295 3590 315
rect 4050 295 4070 315
rect 4230 295 4250 315
rect -145 -95 -125 -75
rect 515 -95 535 -75
rect 1175 -95 1195 -75
rect 1835 -95 1855 -75
rect 2495 -95 2515 -75
rect 3155 -95 3175 -75
rect 3815 -95 3835 -75
<< locali >>
rect 325 800 370 810
rect 325 790 330 800
rect -210 780 330 790
rect 365 790 370 800
rect 985 800 1030 810
rect 985 790 990 800
rect 365 780 990 790
rect 1025 790 1030 800
rect 1645 800 1690 810
rect 1645 790 1650 800
rect 1025 780 1650 790
rect 1685 790 1690 800
rect 2305 800 2350 810
rect 2305 790 2310 800
rect 1685 780 2310 790
rect 2345 790 2350 800
rect 2965 800 3010 810
rect 2965 790 2970 800
rect 2345 780 2970 790
rect 3005 790 3010 800
rect 3625 800 3670 810
rect 3625 790 3630 800
rect 3005 780 3630 790
rect 3665 790 3670 800
rect 3665 780 4330 790
rect -210 770 4330 780
rect -210 730 3800 750
rect -180 650 -160 730
rect -135 700 -95 710
rect -135 680 -125 700
rect -105 690 -95 700
rect 275 700 315 710
rect -105 680 0 690
rect -135 670 0 680
rect -20 650 0 670
rect 275 660 285 700
rect 305 660 315 700
rect -180 640 -140 650
rect -180 355 -170 640
rect -150 355 -140 640
rect -180 345 -140 355
rect -100 640 -60 650
rect -100 355 -90 640
rect -70 355 -60 640
rect -100 345 -60 355
rect -20 640 20 650
rect -20 355 -10 640
rect 10 355 20 640
rect -20 345 20 355
rect 60 640 150 650
rect 60 355 70 640
rect 90 355 120 640
rect 140 355 150 640
rect 275 645 315 660
rect 480 650 500 730
rect 525 700 565 710
rect 525 680 535 700
rect 555 690 565 700
rect 935 700 975 710
rect 555 680 660 690
rect 525 670 660 680
rect 640 650 660 670
rect 935 660 945 700
rect 965 660 975 700
rect 275 495 295 645
rect 480 640 520 650
rect 330 565 370 580
rect 330 525 340 565
rect 360 525 370 565
rect 330 515 370 525
rect 275 485 315 495
rect 275 375 285 485
rect 305 375 315 485
rect 275 365 315 375
rect 375 485 415 495
rect 375 375 385 485
rect 405 375 415 485
rect 375 365 415 375
rect 60 345 150 355
rect -180 320 -160 345
rect -100 320 -80 345
rect -200 300 -160 320
rect -120 310 -75 320
rect -200 265 -180 300
rect -120 290 -115 310
rect -80 290 -75 310
rect -20 305 0 345
rect 395 330 415 365
rect 80 315 120 325
rect 260 320 300 325
rect 80 305 90 315
rect -120 280 -75 290
rect -40 295 90 305
rect 110 295 120 315
rect -40 285 120 295
rect 140 315 300 320
rect 140 300 270 315
rect -200 255 -160 265
rect -200 -30 -190 255
rect -170 -30 -160 255
rect -200 -40 -160 -30
rect -120 255 -80 280
rect -120 -30 -110 255
rect -90 -30 -80 255
rect -120 -40 -80 -30
rect -40 265 -20 285
rect 140 265 160 300
rect 260 295 270 300
rect 290 295 300 315
rect 260 285 300 295
rect 380 310 415 330
rect 480 355 490 640
rect 510 355 520 640
rect 480 345 520 355
rect 560 640 600 650
rect 560 355 570 640
rect 590 355 600 640
rect 560 345 600 355
rect 640 640 680 650
rect 640 355 650 640
rect 670 355 680 640
rect 640 345 680 355
rect 720 640 810 650
rect 720 355 730 640
rect 750 355 780 640
rect 800 355 810 640
rect 935 645 975 660
rect 1140 650 1160 730
rect 1185 700 1225 710
rect 1185 680 1195 700
rect 1215 690 1225 700
rect 1595 700 1635 710
rect 1215 680 1320 690
rect 1185 670 1320 680
rect 1300 650 1320 670
rect 1595 660 1605 700
rect 1625 660 1635 700
rect 935 495 955 645
rect 1140 640 1180 650
rect 990 565 1030 580
rect 990 525 1000 565
rect 1020 525 1030 565
rect 990 515 1030 525
rect 935 485 975 495
rect 935 375 945 485
rect 965 375 975 485
rect 935 365 975 375
rect 1035 485 1075 495
rect 1035 375 1045 485
rect 1065 375 1075 485
rect 1035 365 1075 375
rect 720 345 810 355
rect 480 320 500 345
rect 560 320 580 345
rect 380 265 400 310
rect 460 300 500 320
rect 540 310 585 320
rect 460 265 480 300
rect 540 290 545 310
rect 580 290 585 310
rect 640 305 660 345
rect 1055 330 1075 365
rect 740 315 780 325
rect 920 320 960 325
rect 740 305 750 315
rect 540 280 585 290
rect 620 295 750 305
rect 770 295 780 315
rect 620 285 780 295
rect 800 315 960 320
rect 800 300 930 315
rect -40 255 0 265
rect -40 -30 -30 255
rect -10 -30 0 255
rect -40 -40 0 -30
rect 40 255 80 265
rect 40 -30 50 255
rect 70 -30 80 255
rect 40 -40 80 -30
rect 120 255 160 265
rect 120 -30 130 255
rect 150 -30 160 255
rect 120 -40 160 -30
rect 200 255 240 265
rect 200 -30 210 255
rect 230 -30 240 255
rect 280 255 320 265
rect 280 145 290 255
rect 310 145 320 255
rect 280 135 320 145
rect 380 255 420 265
rect 380 145 390 255
rect 410 145 420 255
rect 380 135 420 145
rect 460 255 500 265
rect 200 -40 240 -30
rect 460 -30 470 255
rect 490 -30 500 255
rect 460 -40 500 -30
rect 540 255 580 280
rect 540 -30 550 255
rect 570 -30 580 255
rect 540 -40 580 -30
rect 620 265 640 285
rect 800 265 820 300
rect 920 295 930 300
rect 950 295 960 315
rect 920 285 960 295
rect 1040 310 1075 330
rect 1140 355 1150 640
rect 1170 355 1180 640
rect 1140 345 1180 355
rect 1220 640 1260 650
rect 1220 355 1230 640
rect 1250 355 1260 640
rect 1220 345 1260 355
rect 1300 640 1340 650
rect 1300 355 1310 640
rect 1330 355 1340 640
rect 1300 345 1340 355
rect 1380 640 1470 650
rect 1380 355 1390 640
rect 1410 355 1440 640
rect 1460 355 1470 640
rect 1595 645 1635 660
rect 1800 650 1820 730
rect 1845 700 1885 710
rect 1845 680 1855 700
rect 1875 690 1885 700
rect 2255 700 2295 710
rect 1875 680 1980 690
rect 1845 670 1980 680
rect 1960 650 1980 670
rect 2255 660 2265 700
rect 2285 660 2295 700
rect 1595 495 1615 645
rect 1800 640 1840 650
rect 1650 565 1690 580
rect 1650 525 1660 565
rect 1680 525 1690 565
rect 1650 515 1690 525
rect 1595 485 1635 495
rect 1595 375 1605 485
rect 1625 375 1635 485
rect 1595 365 1635 375
rect 1695 485 1735 495
rect 1695 375 1705 485
rect 1725 375 1735 485
rect 1695 365 1735 375
rect 1380 345 1470 355
rect 1140 320 1160 345
rect 1220 320 1240 345
rect 1040 265 1060 310
rect 1120 300 1160 320
rect 1200 310 1245 320
rect 1120 265 1140 300
rect 1200 290 1205 310
rect 1240 290 1245 310
rect 1300 305 1320 345
rect 1715 330 1735 365
rect 1400 315 1440 325
rect 1580 320 1620 325
rect 1400 305 1410 315
rect 1200 280 1245 290
rect 1280 295 1410 305
rect 1430 295 1440 315
rect 1280 285 1440 295
rect 1460 315 1620 320
rect 1460 300 1590 315
rect 620 255 660 265
rect 620 -30 630 255
rect 650 -30 660 255
rect 620 -40 660 -30
rect 700 255 740 265
rect 700 -30 710 255
rect 730 -30 740 255
rect 700 -40 740 -30
rect 780 255 820 265
rect 780 -30 790 255
rect 810 -30 820 255
rect 780 -40 820 -30
rect 860 255 900 265
rect 860 -30 870 255
rect 890 -30 900 255
rect 940 255 980 265
rect 940 145 950 255
rect 970 145 980 255
rect 940 135 980 145
rect 1040 255 1080 265
rect 1040 145 1050 255
rect 1070 145 1080 255
rect 1040 135 1080 145
rect 1120 255 1160 265
rect 860 -40 900 -30
rect 1120 -30 1130 255
rect 1150 -30 1160 255
rect 1120 -40 1160 -30
rect 1200 255 1240 280
rect 1200 -30 1210 255
rect 1230 -30 1240 255
rect 1200 -40 1240 -30
rect 1280 265 1300 285
rect 1460 265 1480 300
rect 1580 295 1590 300
rect 1610 295 1620 315
rect 1580 285 1620 295
rect 1700 310 1735 330
rect 1800 355 1810 640
rect 1830 355 1840 640
rect 1800 345 1840 355
rect 1880 640 1920 650
rect 1880 355 1890 640
rect 1910 355 1920 640
rect 1880 345 1920 355
rect 1960 640 2000 650
rect 1960 355 1970 640
rect 1990 355 2000 640
rect 1960 345 2000 355
rect 2040 640 2130 650
rect 2040 355 2050 640
rect 2070 355 2100 640
rect 2120 355 2130 640
rect 2255 645 2295 660
rect 2460 650 2480 730
rect 2505 700 2545 710
rect 2505 680 2515 700
rect 2535 690 2545 700
rect 2915 700 2955 710
rect 2535 680 2640 690
rect 2505 670 2640 680
rect 2620 650 2640 670
rect 2915 660 2925 700
rect 2945 660 2955 700
rect 2255 495 2275 645
rect 2460 640 2500 650
rect 2310 565 2350 580
rect 2310 525 2320 565
rect 2340 525 2350 565
rect 2310 515 2350 525
rect 2255 485 2295 495
rect 2255 375 2265 485
rect 2285 375 2295 485
rect 2255 365 2295 375
rect 2355 485 2395 495
rect 2355 375 2365 485
rect 2385 375 2395 485
rect 2355 365 2395 375
rect 2040 345 2130 355
rect 1800 320 1820 345
rect 1880 320 1900 345
rect 1700 265 1720 310
rect 1780 300 1820 320
rect 1860 310 1905 320
rect 1780 265 1800 300
rect 1860 290 1865 310
rect 1900 290 1905 310
rect 1960 305 1980 345
rect 2375 330 2395 365
rect 2060 315 2100 325
rect 2240 320 2280 325
rect 2060 305 2070 315
rect 1860 280 1905 290
rect 1940 295 2070 305
rect 2090 295 2100 315
rect 1940 285 2100 295
rect 2120 315 2280 320
rect 2120 300 2250 315
rect 1280 255 1320 265
rect 1280 -30 1290 255
rect 1310 -30 1320 255
rect 1280 -40 1320 -30
rect 1360 255 1400 265
rect 1360 -30 1370 255
rect 1390 -30 1400 255
rect 1360 -40 1400 -30
rect 1440 255 1480 265
rect 1440 -30 1450 255
rect 1470 -30 1480 255
rect 1440 -40 1480 -30
rect 1520 255 1560 265
rect 1520 -30 1530 255
rect 1550 -30 1560 255
rect 1600 255 1640 265
rect 1600 145 1610 255
rect 1630 145 1640 255
rect 1600 135 1640 145
rect 1700 255 1740 265
rect 1700 145 1710 255
rect 1730 145 1740 255
rect 1700 135 1740 145
rect 1780 255 1820 265
rect 1520 -40 1560 -30
rect 1780 -30 1790 255
rect 1810 -30 1820 255
rect 1780 -40 1820 -30
rect 1860 255 1900 280
rect 1860 -30 1870 255
rect 1890 -30 1900 255
rect 1860 -40 1900 -30
rect 1940 265 1960 285
rect 2120 265 2140 300
rect 2240 295 2250 300
rect 2270 295 2280 315
rect 2240 285 2280 295
rect 2360 310 2395 330
rect 2460 355 2470 640
rect 2490 355 2500 640
rect 2460 345 2500 355
rect 2540 640 2580 650
rect 2540 355 2550 640
rect 2570 355 2580 640
rect 2540 345 2580 355
rect 2620 640 2660 650
rect 2620 355 2630 640
rect 2650 355 2660 640
rect 2620 345 2660 355
rect 2700 640 2790 650
rect 2700 355 2710 640
rect 2730 355 2760 640
rect 2780 355 2790 640
rect 2915 645 2955 660
rect 3120 650 3140 730
rect 3165 700 3205 710
rect 3165 680 3175 700
rect 3195 690 3205 700
rect 3575 700 3615 710
rect 3195 680 3300 690
rect 3165 670 3300 680
rect 3280 650 3300 670
rect 3575 660 3585 700
rect 3605 660 3615 700
rect 2915 495 2935 645
rect 3120 640 3160 650
rect 2970 565 3010 580
rect 2970 525 2980 565
rect 3000 525 3010 565
rect 2970 515 3010 525
rect 2915 485 2955 495
rect 2915 375 2925 485
rect 2945 375 2955 485
rect 2915 365 2955 375
rect 3015 485 3055 495
rect 3015 375 3025 485
rect 3045 375 3055 485
rect 3015 365 3055 375
rect 2700 345 2790 355
rect 2460 320 2480 345
rect 2540 320 2560 345
rect 2360 265 2380 310
rect 2440 300 2480 320
rect 2520 310 2565 320
rect 2440 265 2460 300
rect 2520 290 2525 310
rect 2560 290 2565 310
rect 2620 305 2640 345
rect 3035 330 3055 365
rect 2720 315 2760 325
rect 2900 320 2940 325
rect 2720 305 2730 315
rect 2520 280 2565 290
rect 2600 295 2730 305
rect 2750 295 2760 315
rect 2600 285 2760 295
rect 2780 315 2940 320
rect 2780 300 2910 315
rect 1940 255 1980 265
rect 1940 -30 1950 255
rect 1970 -30 1980 255
rect 1940 -40 1980 -30
rect 2020 255 2060 265
rect 2020 -30 2030 255
rect 2050 -30 2060 255
rect 2020 -40 2060 -30
rect 2100 255 2140 265
rect 2100 -30 2110 255
rect 2130 -30 2140 255
rect 2100 -40 2140 -30
rect 2180 255 2220 265
rect 2180 -30 2190 255
rect 2210 -30 2220 255
rect 2260 255 2300 265
rect 2260 145 2270 255
rect 2290 145 2300 255
rect 2260 135 2300 145
rect 2360 255 2400 265
rect 2360 145 2370 255
rect 2390 145 2400 255
rect 2360 135 2400 145
rect 2440 255 2480 265
rect 2180 -40 2220 -30
rect 2440 -30 2450 255
rect 2470 -30 2480 255
rect 2440 -40 2480 -30
rect 2520 255 2560 280
rect 2520 -30 2530 255
rect 2550 -30 2560 255
rect 2520 -40 2560 -30
rect 2600 265 2620 285
rect 2780 265 2800 300
rect 2900 295 2910 300
rect 2930 295 2940 315
rect 2900 285 2940 295
rect 3020 310 3055 330
rect 3120 355 3130 640
rect 3150 355 3160 640
rect 3120 345 3160 355
rect 3200 640 3240 650
rect 3200 355 3210 640
rect 3230 355 3240 640
rect 3200 345 3240 355
rect 3280 640 3320 650
rect 3280 355 3290 640
rect 3310 355 3320 640
rect 3280 345 3320 355
rect 3360 640 3450 650
rect 3360 355 3370 640
rect 3390 355 3420 640
rect 3440 355 3450 640
rect 3575 645 3615 660
rect 3780 650 3800 730
rect 3825 700 3865 710
rect 3825 680 3835 700
rect 3855 690 3865 700
rect 4235 700 4275 710
rect 3855 680 3960 690
rect 3825 670 3960 680
rect 3940 650 3960 670
rect 4235 660 4245 700
rect 4265 660 4275 700
rect 3575 495 3595 645
rect 3780 640 3820 650
rect 3630 565 3670 580
rect 3630 525 3640 565
rect 3660 525 3670 565
rect 3630 515 3670 525
rect 3575 485 3615 495
rect 3575 375 3585 485
rect 3605 375 3615 485
rect 3575 365 3615 375
rect 3675 485 3715 495
rect 3675 375 3685 485
rect 3705 375 3715 485
rect 3675 365 3715 375
rect 3360 345 3450 355
rect 3120 320 3140 345
rect 3200 320 3220 345
rect 3020 265 3040 310
rect 3100 300 3140 320
rect 3180 310 3225 320
rect 3100 265 3120 300
rect 3180 290 3185 310
rect 3220 290 3225 310
rect 3280 305 3300 345
rect 3695 330 3715 365
rect 3380 315 3420 325
rect 3560 320 3600 325
rect 3380 305 3390 315
rect 3180 280 3225 290
rect 3260 295 3390 305
rect 3410 295 3420 315
rect 3260 285 3420 295
rect 3440 315 3600 320
rect 3440 300 3570 315
rect 2600 255 2640 265
rect 2600 -30 2610 255
rect 2630 -30 2640 255
rect 2600 -40 2640 -30
rect 2680 255 2720 265
rect 2680 -30 2690 255
rect 2710 -30 2720 255
rect 2680 -40 2720 -30
rect 2760 255 2800 265
rect 2760 -30 2770 255
rect 2790 -30 2800 255
rect 2760 -40 2800 -30
rect 2840 255 2880 265
rect 2840 -30 2850 255
rect 2870 -30 2880 255
rect 2920 255 2960 265
rect 2920 145 2930 255
rect 2950 145 2960 255
rect 2920 135 2960 145
rect 3020 255 3060 265
rect 3020 145 3030 255
rect 3050 145 3060 255
rect 3020 135 3060 145
rect 3100 255 3140 265
rect 2840 -40 2880 -30
rect 3100 -30 3110 255
rect 3130 -30 3140 255
rect 3100 -40 3140 -30
rect 3180 255 3220 280
rect 3180 -30 3190 255
rect 3210 -30 3220 255
rect 3180 -40 3220 -30
rect 3260 265 3280 285
rect 3440 265 3460 300
rect 3560 295 3570 300
rect 3590 295 3600 315
rect 3560 285 3600 295
rect 3680 310 3715 330
rect 3780 355 3790 640
rect 3810 355 3820 640
rect 3780 345 3820 355
rect 3860 640 3900 650
rect 3860 355 3870 640
rect 3890 355 3900 640
rect 3860 345 3900 355
rect 3940 640 3980 650
rect 3940 355 3950 640
rect 3970 355 3980 640
rect 3940 345 3980 355
rect 4020 640 4110 650
rect 4020 355 4030 640
rect 4050 355 4080 640
rect 4100 355 4110 640
rect 4235 645 4275 660
rect 4235 495 4255 645
rect 4310 555 4330 770
rect 4290 545 4330 555
rect 4290 525 4300 545
rect 4320 525 4330 545
rect 4290 515 4330 525
rect 4235 485 4275 495
rect 4235 375 4245 485
rect 4265 375 4275 485
rect 4235 365 4275 375
rect 4335 485 4375 495
rect 4335 375 4345 485
rect 4365 375 4375 485
rect 4335 365 4375 375
rect 4020 345 4110 355
rect 3780 320 3800 345
rect 3860 320 3880 345
rect 3680 265 3700 310
rect 3760 300 3800 320
rect 3840 310 3885 320
rect 3760 265 3780 300
rect 3840 290 3845 310
rect 3880 290 3885 310
rect 3940 305 3960 345
rect 4355 330 4375 365
rect 4040 315 4080 325
rect 4220 320 4260 325
rect 4040 305 4050 315
rect 3840 280 3885 290
rect 3920 295 4050 305
rect 4070 295 4080 315
rect 3920 285 4080 295
rect 4100 315 4260 320
rect 4100 300 4230 315
rect 3260 255 3300 265
rect 3260 -30 3270 255
rect 3290 -30 3300 255
rect 3260 -40 3300 -30
rect 3340 255 3380 265
rect 3340 -30 3350 255
rect 3370 -30 3380 255
rect 3340 -40 3380 -30
rect 3420 255 3460 265
rect 3420 -30 3430 255
rect 3450 -30 3460 255
rect 3420 -40 3460 -30
rect 3500 255 3540 265
rect 3500 -30 3510 255
rect 3530 -30 3540 255
rect 3580 255 3620 265
rect 3580 145 3590 255
rect 3610 145 3620 255
rect 3580 135 3620 145
rect 3680 255 3720 265
rect 3680 145 3690 255
rect 3710 145 3720 255
rect 3680 135 3720 145
rect 3760 255 3800 265
rect 3500 -40 3540 -30
rect 3760 -30 3770 255
rect 3790 -30 3800 255
rect 3760 -40 3800 -30
rect 3840 255 3880 280
rect 3840 -30 3850 255
rect 3870 -30 3880 255
rect 3840 -40 3880 -30
rect 3920 265 3940 285
rect 4100 265 4120 300
rect 4220 295 4230 300
rect 4250 295 4260 315
rect 4220 285 4260 295
rect 4340 310 4375 330
rect 4340 265 4360 310
rect 3920 255 3960 265
rect 3920 -30 3930 255
rect 3950 -30 3960 255
rect 3920 -40 3960 -30
rect 4000 255 4040 265
rect 4000 -30 4010 255
rect 4030 -30 4040 255
rect 4000 -40 4040 -30
rect 4080 255 4120 265
rect 4080 -30 4090 255
rect 4110 -30 4120 255
rect 4080 -40 4120 -30
rect 4160 255 4200 265
rect 4160 -30 4170 255
rect 4190 -30 4200 255
rect 4240 255 4280 265
rect 4240 145 4250 255
rect 4270 145 4280 255
rect 4240 135 4280 145
rect 4340 255 4380 265
rect 4340 145 4350 255
rect 4370 145 4380 255
rect 4340 135 4380 145
rect 4160 -40 4200 -30
rect -155 -75 -115 -65
rect -155 -95 -145 -75
rect -125 -95 -115 -75
rect -155 -105 -115 -95
rect 505 -75 545 -65
rect 505 -95 515 -75
rect 535 -95 545 -75
rect 505 -105 545 -95
rect 1165 -75 1205 -65
rect 1165 -95 1175 -75
rect 1195 -95 1205 -75
rect 1165 -105 1205 -95
rect 1825 -75 1865 -65
rect 1825 -95 1835 -75
rect 1855 -95 1865 -75
rect 1825 -105 1865 -95
rect 2485 -75 2525 -65
rect 2485 -95 2495 -75
rect 2515 -95 2525 -75
rect 2485 -105 2525 -95
rect 3145 -75 3185 -65
rect 3145 -95 3155 -75
rect 3175 -95 3185 -75
rect 3145 -105 3185 -95
rect 3805 -75 3845 -65
rect 3805 -95 3815 -75
rect 3835 -95 3845 -75
rect 3805 -105 3845 -95
<< viali >>
rect 330 780 365 800
rect 990 780 1025 800
rect 1650 780 1685 800
rect 2310 780 2345 800
rect 2970 780 3005 800
rect 3630 780 3665 800
rect 285 660 305 700
rect 70 355 90 640
rect 120 355 140 640
rect 945 660 965 700
rect 340 545 360 565
rect 340 525 360 545
rect -115 290 -80 310
rect 730 355 750 640
rect 780 355 800 640
rect 1605 660 1625 700
rect 1000 545 1020 565
rect 1000 525 1020 545
rect 545 290 580 310
rect 50 -30 70 255
rect 130 220 150 255
rect 210 -30 230 255
rect 290 145 310 255
rect 1390 355 1410 640
rect 1440 355 1460 640
rect 2265 660 2285 700
rect 1660 545 1680 565
rect 1660 525 1680 545
rect 1205 290 1240 310
rect 710 -30 730 255
rect 790 220 810 255
rect 870 -30 890 255
rect 950 145 970 255
rect 2050 355 2070 640
rect 2100 355 2120 640
rect 2925 660 2945 700
rect 2320 545 2340 565
rect 2320 525 2340 545
rect 1865 290 1900 310
rect 1370 -30 1390 255
rect 1450 220 1470 255
rect 1530 -30 1550 255
rect 1610 145 1630 255
rect 2710 355 2730 640
rect 2760 355 2780 640
rect 3585 660 3605 700
rect 2980 545 3000 565
rect 2980 525 3000 545
rect 2525 290 2560 310
rect 2030 -30 2050 255
rect 2110 220 2130 255
rect 2190 -30 2210 255
rect 2270 145 2290 255
rect 3370 355 3390 640
rect 3420 355 3440 640
rect 4245 660 4265 700
rect 3640 545 3660 565
rect 3640 525 3660 545
rect 3185 290 3220 310
rect 2690 -30 2710 255
rect 2770 220 2790 255
rect 2850 -30 2870 255
rect 2930 145 2950 255
rect 4030 355 4050 640
rect 4080 355 4100 640
rect 3845 290 3880 310
rect 3350 -30 3370 255
rect 3430 220 3450 255
rect 3510 -30 3530 255
rect 3590 145 3610 255
rect 4010 -30 4030 255
rect 4090 220 4110 255
rect 4170 -30 4190 255
rect 4250 145 4270 255
<< metal1 >>
rect 275 710 295 820
rect 325 800 370 810
rect 325 780 330 800
rect 365 780 370 800
rect 325 770 370 780
rect 275 700 315 710
rect 275 660 285 700
rect 305 660 315 700
rect 60 640 150 650
rect 275 645 315 660
rect 60 440 70 640
rect -205 355 70 440
rect 90 355 120 640
rect 140 440 150 640
rect 330 565 370 770
rect 935 710 955 820
rect 985 800 1030 810
rect 985 780 990 800
rect 1025 780 1030 800
rect 985 770 1030 780
rect 935 700 975 710
rect 935 660 945 700
rect 965 660 975 700
rect 330 525 340 565
rect 360 525 370 565
rect 330 515 370 525
rect 720 640 810 650
rect 935 645 975 660
rect 720 440 730 640
rect 140 355 730 440
rect 750 355 780 640
rect 800 440 810 640
rect 990 565 1030 770
rect 1595 710 1615 820
rect 1645 800 1690 810
rect 1645 780 1650 800
rect 1685 780 1690 800
rect 1645 770 1690 780
rect 1595 700 1635 710
rect 1595 660 1605 700
rect 1625 660 1635 700
rect 990 525 1000 565
rect 1020 525 1030 565
rect 990 515 1030 525
rect 1380 640 1470 650
rect 1595 645 1635 660
rect 1380 440 1390 640
rect 800 355 1390 440
rect 1410 355 1440 640
rect 1460 440 1470 640
rect 1650 565 1690 770
rect 2255 710 2275 820
rect 2305 800 2350 810
rect 2305 780 2310 800
rect 2345 780 2350 800
rect 2305 770 2350 780
rect 2255 700 2295 710
rect 2255 660 2265 700
rect 2285 660 2295 700
rect 1650 525 1660 565
rect 1680 525 1690 565
rect 1650 515 1690 525
rect 2040 640 2130 650
rect 2255 645 2295 660
rect 2040 440 2050 640
rect 1460 355 2050 440
rect 2070 355 2100 640
rect 2120 440 2130 640
rect 2310 565 2350 770
rect 2915 710 2935 820
rect 2965 800 3010 810
rect 2965 780 2970 800
rect 3005 780 3010 800
rect 2965 770 3010 780
rect 2915 700 2955 710
rect 2915 660 2925 700
rect 2945 660 2955 700
rect 2310 525 2320 565
rect 2340 525 2350 565
rect 2310 515 2350 525
rect 2700 640 2790 650
rect 2915 645 2955 660
rect 2700 440 2710 640
rect 2120 355 2710 440
rect 2730 355 2760 640
rect 2780 440 2790 640
rect 2970 565 3010 770
rect 3575 710 3595 820
rect 3625 800 3670 810
rect 3625 780 3630 800
rect 3665 780 3670 800
rect 3625 770 3670 780
rect 3575 700 3615 710
rect 3575 660 3585 700
rect 3605 660 3615 700
rect 2970 525 2980 565
rect 3000 525 3010 565
rect 2970 515 3010 525
rect 3360 640 3450 650
rect 3575 645 3615 660
rect 3360 440 3370 640
rect 2780 355 3370 440
rect 3390 355 3420 640
rect 3440 440 3450 640
rect 3630 565 3670 770
rect 4235 710 4255 820
rect 4235 700 4275 710
rect 4235 660 4245 700
rect 4265 660 4275 700
rect 3630 525 3640 565
rect 3660 525 3670 565
rect 3630 515 3670 525
rect 4020 640 4110 650
rect 4235 645 4275 660
rect 4020 440 4030 640
rect 3440 355 4030 440
rect 4050 355 4080 640
rect 4100 355 4110 640
rect -205 345 4110 355
rect -120 310 -75 320
rect -120 290 -115 310
rect -80 295 -75 310
rect 540 310 585 320
rect -80 290 160 295
rect -120 280 160 290
rect 540 290 545 310
rect 580 295 585 310
rect 1200 310 1245 320
rect 580 290 820 295
rect 540 280 820 290
rect 1200 290 1205 310
rect 1240 295 1245 310
rect 1860 310 1905 320
rect 1240 290 1480 295
rect 1200 280 1480 290
rect 1860 290 1865 310
rect 1900 295 1905 310
rect 2520 310 2565 320
rect 1900 290 2140 295
rect 1860 280 2140 290
rect 2520 290 2525 310
rect 2560 295 2565 310
rect 3180 310 3225 320
rect 2560 290 2800 295
rect 2520 280 2800 290
rect 3180 290 3185 310
rect 3220 295 3225 310
rect 3840 310 3885 320
rect 3220 290 3460 295
rect 3180 280 3460 290
rect 3840 290 3845 310
rect 3880 295 3885 310
rect 3880 290 4120 295
rect 3840 280 4120 290
rect -205 255 80 265
rect -205 -30 50 255
rect 70 185 80 255
rect 120 255 160 280
rect 120 220 130 255
rect 150 220 160 255
rect 120 210 160 220
rect 200 255 740 265
rect 200 185 210 255
rect 70 -30 210 185
rect 230 145 290 255
rect 310 145 710 255
rect 230 135 710 145
rect 230 -30 240 135
rect -205 -40 240 -30
rect 455 -30 710 135
rect 730 185 740 255
rect 780 255 820 280
rect 780 220 790 255
rect 810 220 820 255
rect 780 210 820 220
rect 860 255 1400 265
rect 860 185 870 255
rect 730 -30 870 185
rect 890 145 950 255
rect 970 145 1370 255
rect 890 135 1370 145
rect 890 -30 900 135
rect 455 -40 900 -30
rect 1115 -30 1370 135
rect 1390 185 1400 255
rect 1440 255 1480 280
rect 1440 220 1450 255
rect 1470 220 1480 255
rect 1440 210 1480 220
rect 1520 255 2060 265
rect 1520 185 1530 255
rect 1390 -30 1530 185
rect 1550 145 1610 255
rect 1630 145 2030 255
rect 1550 135 2030 145
rect 1550 -30 1560 135
rect 1115 -40 1560 -30
rect 1775 -30 2030 135
rect 2050 185 2060 255
rect 2100 255 2140 280
rect 2100 220 2110 255
rect 2130 220 2140 255
rect 2100 210 2140 220
rect 2180 255 2720 265
rect 2180 185 2190 255
rect 2050 -30 2190 185
rect 2210 145 2270 255
rect 2290 145 2690 255
rect 2210 135 2690 145
rect 2210 -30 2220 135
rect 1775 -40 2220 -30
rect 2435 -30 2690 135
rect 2710 185 2720 255
rect 2760 255 2800 280
rect 2760 220 2770 255
rect 2790 220 2800 255
rect 2760 210 2800 220
rect 2840 255 3380 265
rect 2840 185 2850 255
rect 2710 -30 2850 185
rect 2870 145 2930 255
rect 2950 145 3350 255
rect 2870 135 3350 145
rect 2870 -30 2880 135
rect 2435 -40 2880 -30
rect 3095 -30 3350 135
rect 3370 185 3380 255
rect 3420 255 3460 280
rect 3420 220 3430 255
rect 3450 220 3460 255
rect 3420 210 3460 220
rect 3500 255 4040 265
rect 3500 185 3510 255
rect 3370 -30 3510 185
rect 3530 145 3590 255
rect 3610 145 4010 255
rect 3530 135 4010 145
rect 3530 -30 3540 135
rect 3095 -40 3540 -30
rect 3755 -30 4010 135
rect 4030 185 4040 255
rect 4080 255 4120 280
rect 4080 220 4090 255
rect 4110 220 4120 255
rect 4080 210 4120 220
rect 4160 255 4280 265
rect 4160 185 4170 255
rect 4030 -30 4170 185
rect 4190 145 4250 255
rect 4270 145 4280 255
rect 4190 135 4280 145
rect 4190 -30 4200 135
rect 3755 -40 4200 -30
rect 200 -45 240 -40
rect 860 -45 900 -40
rect 1520 -45 1560 -40
rect 2180 -45 2220 -40
rect 2840 -45 2880 -40
rect 3500 -45 3540 -40
rect 4160 -45 4200 -40
<< labels >>
rlabel metal1 -205 390 -205 390 7 VP
rlabel metal1 -205 110 -205 110 7 VN
rlabel locali -135 -105 -135 -105 5 b0in
rlabel locali 525 -105 525 -105 5 b1in
rlabel locali 1185 -105 1185 -105 5 b2in
rlabel locali 1845 -105 1845 -105 5 b3in
rlabel locali 2505 -105 2505 -105 5 b4in
rlabel locali 3165 -105 3165 -105 5 b5in
rlabel locali 3825 -105 3825 -105 5 b6in
rlabel locali -210 740 -210 740 7 Vbn
rlabel locali -210 780 -210 780 7 Vc
rlabel metal1 285 820 285 820 1 branch0
rlabel metal1 945 820 945 820 1 branch1
rlabel metal1 1605 820 1605 820 1 branch2
rlabel metal1 2265 820 2265 820 1 branch3
rlabel metal1 2925 820 2925 820 1 branch4
rlabel metal1 3585 820 3585 820 1 branch5
rlabel metal1 4245 820 4245 820 1 branch6
<< end >>
